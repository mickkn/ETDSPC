-- SOPC_Video.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.03.31.14:42:21

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SOPC_Video is
	port (
		VGA_CLK_from_the_VGA_Controller                     : out   std_logic;                                        --   VGA_Controller_external_interface.CLK
		VGA_HS_from_the_VGA_Controller                      : out   std_logic;                                        --                                    .HS
		VGA_VS_from_the_VGA_Controller                      : out   std_logic;                                        --                                    .VS
		VGA_BLANK_from_the_VGA_Controller                   : out   std_logic;                                        --                                    .BLANK
		VGA_SYNC_from_the_VGA_Controller                    : out   std_logic;                                        --                                    .SYNC
		VGA_R_from_the_VGA_Controller                       : out   std_logic_vector(9 downto 0);                     --                                    .R
		VGA_G_from_the_VGA_Controller                       : out   std_logic_vector(9 downto 0);                     --                                    .G
		VGA_B_from_the_VGA_Controller                       : out   std_logic_vector(9 downto 0);                     --                                    .B
		clk_0                                               : in    std_logic                     := '0';             --                        clk_0_clk_in.clk
		reset_n                                             : in    std_logic                     := '0';             --                  clk_0_clk_in_reset.reset_n
		I2C_SDAT_to_and_from_the_AV_Config                  : inout std_logic                     := '0';             --        AV_Config_external_interface.SDAT
		I2C_SCLK_from_the_AV_Config                         : out   std_logic;                                        --                                    .SCLK
		SRAM_DQ_to_and_from_the_Pixel_Buffer                : inout std_logic_vector(15 downto 0) := (others => '0'); --     Pixel_Buffer_external_interface.DQ
		SRAM_ADDR_from_the_Pixel_Buffer                     : out   std_logic_vector(17 downto 0);                    --                                    .ADDR
		SRAM_LB_N_from_the_Pixel_Buffer                     : out   std_logic;                                        --                                    .LB_N
		SRAM_UB_N_from_the_Pixel_Buffer                     : out   std_logic;                                        --                                    .UB_N
		SRAM_CE_N_from_the_Pixel_Buffer                     : out   std_logic;                                        --                                    .CE_N
		SRAM_OE_N_from_the_Pixel_Buffer                     : out   std_logic;                                        --                                    .OE_N
		SRAM_WE_N_from_the_Pixel_Buffer                     : out   std_logic;                                        --                                    .WE_N
		Video_In_Decoder_external_interface_PIXEL_CLK       : in    std_logic                     := '0';             -- Video_In_Decoder_external_interface.PIXEL_CLK
		Video_In_Decoder_external_interface_LINE_VALID      : in    std_logic                     := '0';             --                                    .LINE_VALID
		Video_In_Decoder_external_interface_FRAME_VALID     : in    std_logic                     := '0';             --                                    .FRAME_VALID
		Video_In_Decoder_external_interface_pixel_clk_reset : in    std_logic                     := '0';             --                                    .pixel_clk_reset
		Video_In_Decoder_external_interface_PIXEL_DATA      : in    std_logic_vector(11 downto 0) := (others => '0'); --                                    .PIXEL_DATA
		vga_clk                                             : out   std_logic;                                        --                                 vga.clk
		sdram_wire_addr                                     : out   std_logic_vector(11 downto 0);                    --                          sdram_wire.addr
		sdram_wire_ba                                       : out   std_logic_vector(1 downto 0);                     --                                    .ba
		sdram_wire_cas_n                                    : out   std_logic;                                        --                                    .cas_n
		sdram_wire_cke                                      : out   std_logic;                                        --                                    .cke
		sdram_wire_cs_n                                     : out   std_logic;                                        --                                    .cs_n
		sdram_wire_dq                                       : inout std_logic_vector(15 downto 0) := (others => '0'); --                                    .dq
		sdram_wire_dqm                                      : out   std_logic_vector(1 downto 0);                     --                                    .dqm
		sdram_wire_ras_n                                    : out   std_logic;                                        --                                    .ras_n
		sdram_wire_we_n                                     : out   std_logic;                                        --                                    .we_n
		lcd_ext_RS                                          : out   std_logic;                                        --                             lcd_ext.RS
		lcd_ext_RW                                          : out   std_logic;                                        --                                    .RW
		lcd_ext_data                                        : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                    .data
		lcd_ext_E                                           : out   std_logic;                                        --                                    .E
		red_leds_ext_export                                 : out   std_logic_vector(7 downto 0);                     --                        red_leds_ext.export
		green_leds_ext_export                               : out   std_logic_vector(7 downto 0);                     --                      green_leds_ext.export
		switch_ext_export                                   : in    std_logic_vector(7 downto 0)  := (others => '0'); --                          switch_ext.export
		altera_up_sd_card_b_SD_cmd                          : inout std_logic                     := '0';             --                   altera_up_sd_card.b_SD_cmd
		altera_up_sd_card_b_SD_dat                          : inout std_logic                     := '0';             --                                    .b_SD_dat
		altera_up_sd_card_b_SD_dat3                         : inout std_logic                     := '0';             --                                    .b_SD_dat3
		altera_up_sd_card_o_SD_clock                        : out   std_logic;                                        --                                    .o_SD_clock
		sdram_clk_clk                                       : out   std_logic;                                        --                           sdram_clk.clk
		restart_export                                      : in    std_logic                     := '0';             --                             restart.export
		debug_export                                        : out   std_logic_vector(7 downto 0)                      --                               debug.export
	);
end entity SOPC_Video;

architecture rtl of SOPC_Video is
	component SOPC_Video_Onchip_Memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component SOPC_Video_Onchip_Memory;

	component SOPC_Video_Dual_Clock_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component SOPC_Video_Dual_Clock_FIFO;

	component SOPC_Video_Pixel_Buffer is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component SOPC_Video_Pixel_Buffer;

	component SOPC_Video_Pixel_Buffer_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component SOPC_Video_Pixel_Buffer_DMA;

	component SOPC_Video_Pixel_RGB_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component SOPC_Video_Pixel_RGB_Resampler;

	component SOPC_Video_VGA_Controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(9 downto 0);                     -- export
			VGA_G         : out std_logic_vector(9 downto 0);                     -- export
			VGA_B         : out std_logic_vector(9 downto 0)                      -- export
		);
	end component SOPC_Video_VGA_Controller;

	component SOPC_Video_Video_In_Decoder is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                     -- data
			PIXEL_CLK                : in  std_logic                     := 'X';             -- export
			LINE_VALID               : in  std_logic                     := 'X';             -- export
			FRAME_VALID              : in  std_logic                     := 'X';             -- export
			pixel_clk_reset          : in  std_logic                     := 'X';             -- export
			PIXEL_DATA               : in  std_logic_vector(11 downto 0) := (others => 'X')  -- export
		);
	end component SOPC_Video_Video_In_Decoder;

	component SOPC_Video_Video_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(7 downto 0)                      -- writedata
		);
	end component SOPC_Video_Video_DMA;

	component SOPC_Video_AV_Config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component SOPC_Video_AV_Config;

	component SOPC_Video_CPU is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_multi_done                       : in  std_logic                     := 'X';             -- done
			E_ci_multi_clk_en                     : out std_logic;                                        -- clk_en
			E_ci_multi_start                      : out std_logic;                                        -- start
			E_ci_result                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                                : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                                : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                                : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                                : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                           : out std_logic;                                        -- readra
			D_ci_readrb                           : out std_logic;                                        -- readrb
			D_ci_writerc                          : out std_logic;                                        -- writerc
			E_ci_dataa                            : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                            : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                      : out std_logic;                                        -- clk
			E_ci_multi_reset                      : out std_logic;                                        -- reset
			W_ci_estatus                          : out std_logic;                                        -- estatus
			W_ci_ipending                         : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component SOPC_Video_CPU;

	component SOPC_Video_Clock_Signals is
		port (
			CLOCK_50    : in  std_logic := 'X'; -- clk
			reset       : in  std_logic := 'X'; -- reset
			sys_clk     : out std_logic;        -- clk
			sys_reset_n : out std_logic;        -- reset_n
			SDRAM_CLK   : out std_logic;        -- clk
			VGA_CLK     : out std_logic         -- clk
		);
	end component SOPC_Video_Clock_Signals;

	component SOPC_Video_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component SOPC_Video_jtag_uart_0;

	component SOPC_Video_video_bayer_resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_data          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic                                         -- valid
		);
	end component SOPC_Video_video_bayer_resampler;

	component SOPC_Video_video_clipper_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_data          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic                                         -- valid
		);
	end component SOPC_Video_video_clipper_0;

	component SOPC_Video_video_scaler_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component SOPC_Video_video_scaler_0;

	component SOPC_Video_video_rgb_resampler_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component SOPC_Video_video_rgb_resampler_0;

	component SOPC_Video_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component SOPC_Video_sysid_qsys_0;

	component SOPC_Video_sdram_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component SOPC_Video_sdram_0;

	component SOPC_Video_timer_system is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component SOPC_Video_timer_system;

	component SOPC_Video_lcd is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component SOPC_Video_lcd;

	component SOPC_Video_red_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component SOPC_Video_red_leds;

	component SOPC_Video_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component SOPC_Video_switch;

	component fpoint_wrapper is
		generic (
			useDivider : integer := 0
		);
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			clk_en : in  std_logic                     := 'X';             -- clk_en
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			n      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- n
			reset  : in  std_logic                     := 'X';             -- reset
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component fpoint_wrapper;

	component Altera_UP_SD_Card_Avalon_Interface is
		port (
			i_avalon_chip_select : in    std_logic                     := 'X';             -- chipselect
			i_avalon_address     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			i_avalon_read        : in    std_logic                     := 'X';             -- read
			i_avalon_write       : in    std_logic                     := 'X';             -- write
			i_avalon_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest : out   std_logic;                                        -- waitrequest
			i_clock              : in    std_logic                     := 'X';             -- clk
			i_reset_n            : in    std_logic                     := 'X';             -- reset_n
			b_SD_cmd             : inout std_logic                     := 'X';             -- export
			b_SD_dat             : inout std_logic                     := 'X';             -- export
			b_SD_dat3            : inout std_logic                     := 'X';             -- export
			o_SD_clock           : out   std_logic                                         -- export
		);
	end component Altera_UP_SD_Card_Avalon_Interface;

	component pixel_scan is
		port (
			avs_s1_write             : in  std_logic                    := 'X';             -- write
			avs_s1_read              : in  std_logic                    := 'X';             -- read
			avs_s1_chipselect        : in  std_logic                    := 'X';             -- chipselect
			avs_s1_address           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s1_writedata         : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			avs_s1_readdata          : out std_logic_vector(7 downto 0);                    -- readdata
			ast_sink_ready           : out std_logic;                                       -- ready
			ast_sink_valid           : in  std_logic                    := 'X';             -- valid
			ast_sink_startofpacket   : in  std_logic                    := 'X';             -- startofpacket
			ast_sink_endofpacket     : in  std_logic                    := 'X';             -- endofpacket
			ast_sink_data            : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			clk                      : in  std_logic                    := 'X';             -- clk
			reset_n                  : in  std_logic                    := 'X';             -- reset_n
			avs_s1_clk               : in  std_logic                    := 'X';             -- clk
			avs_s1_reset_n           : in  std_logic                    := 'X';             -- reset_n
			ast_source_valid         : out std_logic;                                       -- valid
			ast_source_endofpacket   : out std_logic;                                       -- endofpacket
			ast_source_data          : out std_logic_vector(7 downto 0);                    -- data
			ast_source_startofpacket : out std_logic;                                       -- startofpacket
			ast_source_ready         : in  std_logic                    := 'X';             -- ready
			debug_state              : out std_logic_vector(7 downto 0);                    -- export
			restart                  : in  std_logic                    := 'X'              -- export
		);
	end component pixel_scan;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result         : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra         : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb         : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc        : in  std_logic                     := 'X';             -- writerc
			ci_slave_a              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus        : in  std_logic                     := 'X';             -- estatus
			ci_slave_multi_clk      : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset    : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken    : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_start    : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done     : out std_logic;                                        -- done
			comb_ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab    : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n        : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra   : out std_logic;                                        -- readra
			comb_ci_master_readrb   : out std_logic;                                        -- readrb
			comb_ci_master_writerc  : out std_logic;                                        -- writerc
			comb_ci_master_a        : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b        : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c        : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus  : out std_logic;                                        -- estatus
			multi_ci_master_clk     : out std_logic;                                        -- clk
			multi_ci_master_reset   : out std_logic;                                        -- reset
			multi_ci_master_clken   : out std_logic;                                        -- clk_en
			multi_ci_master_start   : out std_logic;                                        -- start
			multi_ci_master_done    : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa   : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab   : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n       : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra  : out std_logic;                                        -- readra
			multi_ci_master_readrb  : out std_logic;                                        -- readrb
			multi_ci_master_writerc : out std_logic;                                        -- writerc
			multi_ci_master_a       : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b       : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c       : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_multi_dataa    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result   : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra   : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb   : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc  : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c        : in  std_logic_vector(4 downto 0)  := (others => 'X')  -- multi_c
		);
	end component altera_customins_master_translator;

	component SOPC_Video_CPU_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic;                                        -- done
			ci_master0_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra   : out std_logic;                                        -- readra
			ci_master0_readrb   : out std_logic;                                        -- readrb
			ci_master0_writerc  : out std_logic;                                        -- writerc
			ci_master0_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus  : out std_logic;                                        -- estatus
			ci_master0_clk      : out std_logic;                                        -- clk
			ci_master0_reset    : out std_logic;                                        -- reset
			ci_master0_clken    : out std_logic;                                        -- clk_en
			ci_master0_start    : out std_logic;                                        -- start
			ci_master0_done     : in  std_logic                     := 'X'              -- done
		);
	end component SOPC_Video_CPU_custom_instruction_master_multi_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result    : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra    : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb    : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc   : in  std_logic                     := 'X';             -- writerc
			ci_slave_a         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus   : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk       : in  std_logic                     := 'X';             -- clk
			ci_slave_clken     : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset     : in  std_logic                     := 'X';             -- reset
			ci_slave_start     : in  std_logic                     := 'X';             -- start
			ci_slave_done      : out std_logic;                                        -- done
			ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n        : out std_logic_vector(1 downto 0);                     -- n
			ci_master_clk      : out std_logic;                                        -- clk
			ci_master_clken    : out std_logic;                                        -- clk_en
			ci_master_reset    : out std_logic;                                        -- reset
			ci_master_start    : out std_logic;                                        -- start
			ci_master_done     : in  std_logic                     := 'X';             -- done
			ci_master_readra   : out std_logic;                                        -- readra
			ci_master_readrb   : out std_logic;                                        -- readrb
			ci_master_writerc  : out std_logic;                                        -- writerc
			ci_master_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus  : out std_logic                                         -- estatus
		);
	end component altera_customins_slave_translator;

	component SOPC_Video_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_addr_router;

	component SOPC_Video_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_addr_router_001;

	component SOPC_Video_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_addr_router_002;

	component SOPC_Video_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_id_router;

	component SOPC_Video_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(90 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_id_router_002;

	component SOPC_Video_id_router_003 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(90 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_id_router_003;

	component SOPC_Video_id_router_004 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(108 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_id_router_004;

	component SOPC_Video_id_router_016 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_id_router_016;

	component SOPC_Video_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(108 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(108 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(108 downto 0);                    -- data
			src2_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_demux;

	component SOPC_Video_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			sink_ready          : out std_logic;                                         -- ready
			sink_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready          : in  std_logic                      := 'X';             -- ready
			src0_valid          : out std_logic;                                         -- valid
			src0_data           : out std_logic_vector(108 downto 0);                    -- data
			src0_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket  : out std_logic;                                         -- startofpacket
			src0_endofpacket    : out std_logic;                                         -- endofpacket
			src1_ready          : in  std_logic                      := 'X';             -- ready
			src1_valid          : out std_logic;                                         -- valid
			src1_data           : out std_logic_vector(108 downto 0);                    -- data
			src1_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src1_startofpacket  : out std_logic;                                         -- startofpacket
			src1_endofpacket    : out std_logic;                                         -- endofpacket
			src2_ready          : in  std_logic                      := 'X';             -- ready
			src2_valid          : out std_logic;                                         -- valid
			src2_data           : out std_logic_vector(108 downto 0);                    -- data
			src2_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src2_startofpacket  : out std_logic;                                         -- startofpacket
			src2_endofpacket    : out std_logic;                                         -- endofpacket
			src3_ready          : in  std_logic                      := 'X';             -- ready
			src3_valid          : out std_logic;                                         -- valid
			src3_data           : out std_logic_vector(108 downto 0);                    -- data
			src3_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src3_startofpacket  : out std_logic;                                         -- startofpacket
			src3_endofpacket    : out std_logic;                                         -- endofpacket
			src4_ready          : in  std_logic                      := 'X';             -- ready
			src4_valid          : out std_logic;                                         -- valid
			src4_data           : out std_logic_vector(108 downto 0);                    -- data
			src4_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src4_startofpacket  : out std_logic;                                         -- startofpacket
			src4_endofpacket    : out std_logic;                                         -- endofpacket
			src5_ready          : in  std_logic                      := 'X';             -- ready
			src5_valid          : out std_logic;                                         -- valid
			src5_data           : out std_logic_vector(108 downto 0);                    -- data
			src5_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src5_startofpacket  : out std_logic;                                         -- startofpacket
			src5_endofpacket    : out std_logic;                                         -- endofpacket
			src6_ready          : in  std_logic                      := 'X';             -- ready
			src6_valid          : out std_logic;                                         -- valid
			src6_data           : out std_logic_vector(108 downto 0);                    -- data
			src6_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src6_startofpacket  : out std_logic;                                         -- startofpacket
			src6_endofpacket    : out std_logic;                                         -- endofpacket
			src7_ready          : in  std_logic                      := 'X';             -- ready
			src7_valid          : out std_logic;                                         -- valid
			src7_data           : out std_logic_vector(108 downto 0);                    -- data
			src7_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src7_startofpacket  : out std_logic;                                         -- startofpacket
			src7_endofpacket    : out std_logic;                                         -- endofpacket
			src8_ready          : in  std_logic                      := 'X';             -- ready
			src8_valid          : out std_logic;                                         -- valid
			src8_data           : out std_logic_vector(108 downto 0);                    -- data
			src8_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src8_startofpacket  : out std_logic;                                         -- startofpacket
			src8_endofpacket    : out std_logic;                                         -- endofpacket
			src9_ready          : in  std_logic                      := 'X';             -- ready
			src9_valid          : out std_logic;                                         -- valid
			src9_data           : out std_logic_vector(108 downto 0);                    -- data
			src9_channel        : out std_logic_vector(16 downto 0);                     -- channel
			src9_startofpacket  : out std_logic;                                         -- startofpacket
			src9_endofpacket    : out std_logic;                                         -- endofpacket
			src10_ready         : in  std_logic                      := 'X';             -- ready
			src10_valid         : out std_logic;                                         -- valid
			src10_data          : out std_logic_vector(108 downto 0);                    -- data
			src10_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src10_startofpacket : out std_logic;                                         -- startofpacket
			src10_endofpacket   : out std_logic;                                         -- endofpacket
			src11_ready         : in  std_logic                      := 'X';             -- ready
			src11_valid         : out std_logic;                                         -- valid
			src11_data          : out std_logic_vector(108 downto 0);                    -- data
			src11_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src11_startofpacket : out std_logic;                                         -- startofpacket
			src11_endofpacket   : out std_logic;                                         -- endofpacket
			src12_ready         : in  std_logic                      := 'X';             -- ready
			src12_valid         : out std_logic;                                         -- valid
			src12_data          : out std_logic_vector(108 downto 0);                    -- data
			src12_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src12_startofpacket : out std_logic;                                         -- startofpacket
			src12_endofpacket   : out std_logic;                                         -- endofpacket
			src13_ready         : in  std_logic                      := 'X';             -- ready
			src13_valid         : out std_logic;                                         -- valid
			src13_data          : out std_logic_vector(108 downto 0);                    -- data
			src13_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src13_startofpacket : out std_logic;                                         -- startofpacket
			src13_endofpacket   : out std_logic;                                         -- endofpacket
			src14_ready         : in  std_logic                      := 'X';             -- ready
			src14_valid         : out std_logic;                                         -- valid
			src14_data          : out std_logic_vector(108 downto 0);                    -- data
			src14_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src14_startofpacket : out std_logic;                                         -- startofpacket
			src14_endofpacket   : out std_logic;                                         -- endofpacket
			src15_ready         : in  std_logic                      := 'X';             -- ready
			src15_valid         : out std_logic;                                         -- valid
			src15_data          : out std_logic_vector(108 downto 0);                    -- data
			src15_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src15_startofpacket : out std_logic;                                         -- startofpacket
			src15_endofpacket   : out std_logic;                                         -- endofpacket
			src16_ready         : in  std_logic                      := 'X';             -- ready
			src16_valid         : out std_logic;                                         -- valid
			src16_data          : out std_logic_vector(108 downto 0);                    -- data
			src16_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src16_startofpacket : out std_logic;                                         -- startofpacket
			src16_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_demux_001;

	component SOPC_Video_cmd_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(81 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_demux_002;

	component SOPC_Video_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(108 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_mux;

	component SOPC_Video_cmd_xbar_mux_002 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(90 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_mux_002;

	component SOPC_Video_cmd_xbar_mux_003 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(90 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component SOPC_Video_cmd_xbar_mux_003;

	component SOPC_Video_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(108 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(108 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_demux;

	component SOPC_Video_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(90 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(90 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_demux_002;

	component SOPC_Video_rsp_xbar_demux_003 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(90 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(90 downto 0);                    -- data
			src1_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(90 downto 0);                    -- data
			src2_channel       : out std_logic_vector(16 downto 0);                    -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_demux_003;

	component SOPC_Video_rsp_xbar_demux_004 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(108 downto 0);                    -- data
			src0_channel       : out std_logic_vector(16 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_demux_004;

	component SOPC_Video_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(108 downto 0);                    -- data
			src_channel         : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_mux;

	component SOPC_Video_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_valid            : out std_logic;                                         -- valid
			src_data             : out std_logic_vector(108 downto 0);                    -- data
			src_channel          : out std_logic_vector(16 downto 0);                     -- channel
			src_startofpacket    : out std_logic;                                         -- startofpacket
			src_endofpacket      : out std_logic;                                         -- endofpacket
			sink0_ready          : out std_logic;                                         -- ready
			sink0_valid          : in  std_logic                      := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                         -- ready
			sink1_valid          : in  std_logic                      := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                         -- ready
			sink2_valid          : in  std_logic                      := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                         -- ready
			sink3_valid          : in  std_logic                      := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                         -- ready
			sink4_valid          : in  std_logic                      := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                         -- ready
			sink5_valid          : in  std_logic                      := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                         -- ready
			sink6_valid          : in  std_logic                      := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                         -- ready
			sink7_valid          : in  std_logic                      := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                         -- ready
			sink8_valid          : in  std_logic                      := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                         -- ready
			sink9_valid          : in  std_logic                      := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                         -- ready
			sink10_valid         : in  std_logic                      := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                         -- ready
			sink11_valid         : in  std_logic                      := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                         -- ready
			sink12_valid         : in  std_logic                      := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                         -- ready
			sink13_valid         : in  std_logic                      := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                         -- ready
			sink14_valid         : in  std_logic                      := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                         -- ready
			sink15_valid         : in  std_logic                      := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                         -- ready
			sink16_valid         : in  std_logic                      := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component SOPC_Video_rsp_xbar_mux_001;

	component SOPC_Video_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component SOPC_Video_irq_mapper;

	component sopc_video_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(90 downto 0);                     -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter;

	component sopc_video_width_adapter_003 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(81 downto 0);                     -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter_003;

	component sopc_video_width_adapter_004 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(90 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter_004;

	component sopc_video_width_adapter_006 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(90 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(108 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter_006;

	component sopc_video_width_adapter_009 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(81 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter_009;

	component sopc_video_width_adapter_011 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(81 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(108 downto 0);                    -- data
			out_channel          : out std_logic_vector(16 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_video_width_adapter_011;

	component sopc_video_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(90 downto 0);                    -- data
			source0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component sopc_video_burst_adapter;

	component sopc_video_burst_adapter_002 is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(81 downto 0);                    -- data
			source0_channel       : out std_logic_vector(16 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component sopc_video_burst_adapter_002;

	component sopc_video_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_video_rst_controller;

	component sopc_video_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_video_rst_controller_001;

	component sopc_video_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_video_rst_controller_003;

	component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(109 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(109 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(91 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(91 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(108 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(109 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(109 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(90 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(90 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(91 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(91 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent;

	component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(9 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent;

	component sopc_video_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_video_cpu_instruction_master_translator;

	component sopc_video_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_video_cpu_data_master_translator;

	component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(7 downto 0);                     -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator;

	component sopc_video_video_dma_avalon_dma_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(7 downto 0);                     -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_video_video_dma_avalon_dma_master_translator;

	component sopc_video_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_cpu_jtag_debug_module_translator;

	component sopc_video_onchip_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(11 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_onchip_memory_s1_translator;

	component sopc_video_sdram_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_sdram_0_s1_translator;

	component sopc_video_pixel_buffer_avalon_sram_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(17 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_pixel_buffer_avalon_sram_slave_translator;

	component sopc_video_av_config_avalon_av_config_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_av_config_avalon_av_config_slave_translator;

	component sopc_video_video_dma_avalon_dma_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_video_dma_avalon_dma_control_slave_translator;

	component sopc_video_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_jtag_uart_0_avalon_jtag_slave_translator;

	component sopc_video_sysid_qsys_0_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_sysid_qsys_0_control_slave_translator;

	component sopc_video_timer_system_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_timer_system_s1_translator;

	component sopc_video_lcd_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_lcd_control_slave_translator;

	component sopc_video_red_leds_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_red_leds_s1_translator;

	component sopc_video_switch_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_switch_s1_translator;

	component sopc_video_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator;

	component sopc_video_barcode_scan_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(7 downto 0);                     -- readdata
			uav_writedata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_video_barcode_scan_0_s1_translator;

	component sopc_video_cpu_instruction_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(108 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(108 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component sopc_video_cpu_instruction_master_translator_avalon_universal_master_0_agent;

	component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(7 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(81 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent;

	signal dual_clock_fifo_avalon_dc_buffer_source_endofpacket                                                                           : std_logic;                      -- Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	signal dual_clock_fifo_avalon_dc_buffer_source_valid                                                                                 : std_logic;                      -- Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	signal dual_clock_fifo_avalon_dc_buffer_source_startofpacket                                                                         : std_logic;                      -- Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	signal dual_clock_fifo_avalon_dc_buffer_source_data                                                                                  : std_logic_vector(29 downto 0);  -- Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	signal dual_clock_fifo_avalon_dc_buffer_source_ready                                                                                 : std_logic;                      -- VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	signal clock_signals_sys_clk_clk                                                                                                     : std_logic;                      -- Clock_Signals:sys_clk -> [AV_Config:clk, AV_Config_avalon_av_config_slave_translator:clk, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Altera_UP_SD_Card_Avalon_Interface_0:i_clock, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Barcode_scan_0:avs_s1_clk, Barcode_scan_0:clk, Barcode_scan_0_s1_translator:clk, Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:clk, Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, CPU:clk, CPU_data_master_translator:clk, CPU_data_master_translator_avalon_universal_master_0_agent:clk, CPU_instruction_master_translator:clk, CPU_instruction_master_translator_avalon_universal_master_0_agent:clk, CPU_jtag_debug_module_translator:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Dual_Clock_FIFO:clk_stream_in, Onchip_Memory:clk, Onchip_Memory_s1_translator:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_Buffer:clk, Pixel_Buffer_DMA:clk, Pixel_Buffer_DMA_avalon_control_slave_translator:clk, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:clk, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, Pixel_Buffer_avalon_sram_slave_translator:clk, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_RGB_Resampler:clk, Video_DMA:clk, Video_DMA_avalon_dma_control_slave_translator:clk, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:clk, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Video_DMA_avalon_dma_master_translator:clk, Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, Video_In_Decoder:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, green_leds:clk, green_leds_s1_translator:clk, green_leds_s1_translator_avalon_universal_slave_0_agent:clk, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, lcd:clk, lcd_control_slave_translator:clk, lcd_control_slave_translator_avalon_universal_slave_0_agent:clk, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, red_leds:clk, red_leds_s1_translator:clk, red_leds_s1_translator_avalon_universal_slave_0_agent:clk, red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch:clk, switch_s1_translator:clk, switch_s1_translator_avalon_universal_slave_0_agent:clk, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_system:clk, timer_system_s1_translator:clk, timer_system_s1_translator_avalon_universal_slave_0_agent:clk, timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_timestamp:clk, timer_timestamp_s1_translator:clk, timer_timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_bayer_resampler:clk, video_clipper_0:clk, video_rgb_resampler_0:clk, video_scaler_0:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk]
	signal clock_signals_vga_clk_clk                                                                                                     : std_logic;                      -- Clock_Signals:VGA_CLK -> [vga_clk, Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_001:clk]
	signal pixel_rgb_resampler_avalon_rgb_source_endofpacket                                                                             : std_logic;                      -- Pixel_RGB_Resampler:stream_out_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	signal pixel_rgb_resampler_avalon_rgb_source_valid                                                                                   : std_logic;                      -- Pixel_RGB_Resampler:stream_out_valid -> Dual_Clock_FIFO:stream_in_valid
	signal pixel_rgb_resampler_avalon_rgb_source_startofpacket                                                                           : std_logic;                      -- Pixel_RGB_Resampler:stream_out_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	signal pixel_rgb_resampler_avalon_rgb_source_data                                                                                    : std_logic_vector(29 downto 0);  -- Pixel_RGB_Resampler:stream_out_data -> Dual_Clock_FIFO:stream_in_data
	signal pixel_rgb_resampler_avalon_rgb_source_ready                                                                                   : std_logic;                      -- Dual_Clock_FIFO:stream_in_ready -> Pixel_RGB_Resampler:stream_out_ready
	signal video_in_decoder_avalon_decoder_source_endofpacket                                                                            : std_logic;                      -- Video_In_Decoder:stream_out_endofpacket -> video_bayer_resampler:stream_in_endofpacket
	signal video_in_decoder_avalon_decoder_source_valid                                                                                  : std_logic;                      -- Video_In_Decoder:stream_out_valid -> video_bayer_resampler:stream_in_valid
	signal video_in_decoder_avalon_decoder_source_startofpacket                                                                          : std_logic;                      -- Video_In_Decoder:stream_out_startofpacket -> video_bayer_resampler:stream_in_startofpacket
	signal video_in_decoder_avalon_decoder_source_data                                                                                   : std_logic_vector(7 downto 0);   -- Video_In_Decoder:stream_out_data -> video_bayer_resampler:stream_in_data
	signal video_in_decoder_avalon_decoder_source_ready                                                                                  : std_logic;                      -- video_bayer_resampler:stream_in_ready -> Video_In_Decoder:stream_out_ready
	signal video_bayer_resampler_avalon_bayer_source_endofpacket                                                                         : std_logic;                      -- video_bayer_resampler:stream_out_endofpacket -> video_clipper_0:stream_in_endofpacket
	signal video_bayer_resampler_avalon_bayer_source_valid                                                                               : std_logic;                      -- video_bayer_resampler:stream_out_valid -> video_clipper_0:stream_in_valid
	signal video_bayer_resampler_avalon_bayer_source_startofpacket                                                                       : std_logic;                      -- video_bayer_resampler:stream_out_startofpacket -> video_clipper_0:stream_in_startofpacket
	signal video_bayer_resampler_avalon_bayer_source_data                                                                                : std_logic_vector(23 downto 0);  -- video_bayer_resampler:stream_out_data -> video_clipper_0:stream_in_data
	signal video_bayer_resampler_avalon_bayer_source_ready                                                                               : std_logic;                      -- video_clipper_0:stream_in_ready -> video_bayer_resampler:stream_out_ready
	signal video_rgb_resampler_0_avalon_rgb_source_endofpacket                                                                           : std_logic;                      -- video_rgb_resampler_0:stream_out_endofpacket -> Barcode_scan_0:ast_sink_endofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_valid                                                                                 : std_logic;                      -- video_rgb_resampler_0:stream_out_valid -> Barcode_scan_0:ast_sink_valid
	signal video_rgb_resampler_0_avalon_rgb_source_startofpacket                                                                         : std_logic;                      -- video_rgb_resampler_0:stream_out_startofpacket -> Barcode_scan_0:ast_sink_startofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_data                                                                                  : std_logic_vector(7 downto 0);   -- video_rgb_resampler_0:stream_out_data -> Barcode_scan_0:ast_sink_data
	signal video_rgb_resampler_0_avalon_rgb_source_ready                                                                                 : std_logic;                      -- Barcode_scan_0:ast_sink_ready -> video_rgb_resampler_0:stream_out_ready
	signal pixel_buffer_dma_avalon_pixel_source_endofpacket                                                                              : std_logic;                      -- Pixel_Buffer_DMA:stream_endofpacket -> Pixel_RGB_Resampler:stream_in_endofpacket
	signal pixel_buffer_dma_avalon_pixel_source_valid                                                                                    : std_logic;                      -- Pixel_Buffer_DMA:stream_valid -> Pixel_RGB_Resampler:stream_in_valid
	signal pixel_buffer_dma_avalon_pixel_source_startofpacket                                                                            : std_logic;                      -- Pixel_Buffer_DMA:stream_startofpacket -> Pixel_RGB_Resampler:stream_in_startofpacket
	signal pixel_buffer_dma_avalon_pixel_source_data                                                                                     : std_logic_vector(7 downto 0);   -- Pixel_Buffer_DMA:stream_data -> Pixel_RGB_Resampler:stream_in_data
	signal pixel_buffer_dma_avalon_pixel_source_ready                                                                                    : std_logic;                      -- Pixel_RGB_Resampler:stream_in_ready -> Pixel_Buffer_DMA:stream_ready
	signal video_clipper_0_avalon_clipper_source_endofpacket                                                                             : std_logic;                      -- video_clipper_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	signal video_clipper_0_avalon_clipper_source_valid                                                                                   : std_logic;                      -- video_clipper_0:stream_out_valid -> video_scaler_0:stream_in_valid
	signal video_clipper_0_avalon_clipper_source_startofpacket                                                                           : std_logic;                      -- video_clipper_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	signal video_clipper_0_avalon_clipper_source_data                                                                                    : std_logic_vector(23 downto 0);  -- video_clipper_0:stream_out_data -> video_scaler_0:stream_in_data
	signal video_clipper_0_avalon_clipper_source_ready                                                                                   : std_logic;                      -- video_scaler_0:stream_in_ready -> video_clipper_0:stream_out_ready
	signal video_scaler_0_avalon_scaler_source_endofpacket                                                                               : std_logic;                      -- video_scaler_0:stream_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	signal video_scaler_0_avalon_scaler_source_valid                                                                                     : std_logic;                      -- video_scaler_0:stream_out_valid -> video_rgb_resampler_0:stream_in_valid
	signal video_scaler_0_avalon_scaler_source_startofpacket                                                                             : std_logic;                      -- video_scaler_0:stream_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	signal video_scaler_0_avalon_scaler_source_data                                                                                      : std_logic_vector(23 downto 0);  -- video_scaler_0:stream_out_data -> video_rgb_resampler_0:stream_in_data
	signal video_scaler_0_avalon_scaler_source_ready                                                                                     : std_logic;                      -- video_rgb_resampler_0:stream_in_ready -> video_scaler_0:stream_out_ready
	signal barcode_scan_0_avalon_streaming_source_endofpacket                                                                            : std_logic;                      -- Barcode_scan_0:ast_source_endofpacket -> Video_DMA:stream_endofpacket
	signal barcode_scan_0_avalon_streaming_source_valid                                                                                  : std_logic;                      -- Barcode_scan_0:ast_source_valid -> Video_DMA:stream_valid
	signal barcode_scan_0_avalon_streaming_source_startofpacket                                                                          : std_logic;                      -- Barcode_scan_0:ast_source_startofpacket -> Video_DMA:stream_startofpacket
	signal barcode_scan_0_avalon_streaming_source_data                                                                                   : std_logic_vector(7 downto 0);   -- Barcode_scan_0:ast_source_data -> Video_DMA:stream_data
	signal barcode_scan_0_avalon_streaming_source_ready                                                                                  : std_logic;                      -- Video_DMA:stream_ready -> Barcode_scan_0:ast_source_ready
	signal cpu_custom_instruction_master_result                                                                                          : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_translator:ci_slave_result -> CPU:E_ci_result
	signal cpu_custom_instruction_master_b                                                                                               : std_logic_vector(4 downto 0);   -- CPU:D_ci_b -> CPU_custom_instruction_master_translator:ci_slave_b
	signal cpu_custom_instruction_master_c                                                                                               : std_logic_vector(4 downto 0);   -- CPU:D_ci_c -> CPU_custom_instruction_master_translator:ci_slave_c
	signal cpu_custom_instruction_master_done                                                                                            : std_logic;                      -- CPU_custom_instruction_master_translator:ci_slave_multi_done -> CPU:E_ci_multi_done
	signal cpu_custom_instruction_master_clk_en                                                                                          : std_logic;                      -- CPU:E_ci_multi_clk_en -> CPU_custom_instruction_master_translator:ci_slave_multi_clken
	signal cpu_custom_instruction_master_a                                                                                               : std_logic_vector(4 downto 0);   -- CPU:D_ci_a -> CPU_custom_instruction_master_translator:ci_slave_a
	signal cpu_custom_instruction_master_n                                                                                               : std_logic_vector(7 downto 0);   -- CPU:D_ci_n -> CPU_custom_instruction_master_translator:ci_slave_n
	signal cpu_custom_instruction_master_writerc                                                                                         : std_logic;                      -- CPU:D_ci_writerc -> CPU_custom_instruction_master_translator:ci_slave_writerc
	signal cpu_custom_instruction_master_ipending                                                                                        : std_logic_vector(31 downto 0);  -- CPU:W_ci_ipending -> CPU_custom_instruction_master_translator:ci_slave_ipending
	signal cpu_custom_instruction_master_clk                                                                                             : std_logic;                      -- CPU:E_ci_multi_clock -> CPU_custom_instruction_master_translator:ci_slave_multi_clk
	signal cpu_custom_instruction_master_start                                                                                           : std_logic;                      -- CPU:E_ci_multi_start -> CPU_custom_instruction_master_translator:ci_slave_multi_start
	signal cpu_custom_instruction_master_dataa                                                                                           : std_logic_vector(31 downto 0);  -- CPU:E_ci_dataa -> CPU_custom_instruction_master_translator:ci_slave_dataa
	signal cpu_custom_instruction_master_readra                                                                                          : std_logic;                      -- CPU:D_ci_readra -> CPU_custom_instruction_master_translator:ci_slave_readra
	signal cpu_custom_instruction_master_reset                                                                                           : std_logic;                      -- CPU:E_ci_multi_reset -> CPU_custom_instruction_master_translator:ci_slave_multi_reset
	signal cpu_custom_instruction_master_datab                                                                                           : std_logic_vector(31 downto 0);  -- CPU:E_ci_datab -> CPU_custom_instruction_master_translator:ci_slave_datab
	signal cpu_custom_instruction_master_readrb                                                                                          : std_logic;                      -- CPU:D_ci_readrb -> CPU_custom_instruction_master_translator:ci_slave_readrb
	signal cpu_custom_instruction_master_estatus                                                                                         : std_logic;                      -- CPU:W_ci_estatus -> CPU_custom_instruction_master_translator:ci_slave_estatus
	signal cpu_custom_instruction_master_translator_multi_ci_master_result                                                               : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_xconnect:ci_slave_result -> CPU_custom_instruction_master_translator:multi_ci_master_result
	signal cpu_custom_instruction_master_translator_multi_ci_master_b                                                                    : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_translator:multi_ci_master_b -> CPU_custom_instruction_master_multi_xconnect:ci_slave_b
	signal cpu_custom_instruction_master_translator_multi_ci_master_c                                                                    : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_translator:multi_ci_master_c -> CPU_custom_instruction_master_multi_xconnect:ci_slave_c
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk_en                                                               : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_clken -> CPU_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal cpu_custom_instruction_master_translator_multi_ci_master_done                                                                 : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_slave_done -> CPU_custom_instruction_master_translator:multi_ci_master_done
	signal cpu_custom_instruction_master_translator_multi_ci_master_a                                                                    : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_translator:multi_ci_master_a -> CPU_custom_instruction_master_multi_xconnect:ci_slave_a
	signal cpu_custom_instruction_master_translator_multi_ci_master_n                                                                    : std_logic_vector(7 downto 0);   -- CPU_custom_instruction_master_translator:multi_ci_master_n -> CPU_custom_instruction_master_multi_xconnect:ci_slave_n
	signal cpu_custom_instruction_master_translator_multi_ci_master_writerc                                                              : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_writerc -> CPU_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk                                                                  : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_clk -> CPU_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal cpu_custom_instruction_master_translator_multi_ci_master_start                                                                : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_start -> CPU_custom_instruction_master_multi_xconnect:ci_slave_start
	signal cpu_custom_instruction_master_translator_multi_ci_master_dataa                                                                : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_translator:multi_ci_master_dataa -> CPU_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal cpu_custom_instruction_master_translator_multi_ci_master_readra                                                               : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_readra -> CPU_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal cpu_custom_instruction_master_translator_multi_ci_master_reset                                                                : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_reset -> CPU_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal cpu_custom_instruction_master_translator_multi_ci_master_datab                                                                : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_translator:multi_ci_master_datab -> CPU_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal cpu_custom_instruction_master_translator_multi_ci_master_readrb                                                               : std_logic;                      -- CPU_custom_instruction_master_translator:multi_ci_master_readrb -> CPU_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_result                                                                : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_slave_translator0:ci_slave_result -> CPU_custom_instruction_master_multi_xconnect:ci_master0_result
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_b                                                                     : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_multi_xconnect:ci_master0_b -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_c                                                                     : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_multi_xconnect:ci_master0_c -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_done                                                                  : std_logic;                      -- CPU_custom_instruction_master_multi_slave_translator0:ci_slave_done -> CPU_custom_instruction_master_multi_xconnect:ci_master0_done
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en                                                                : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_clken -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_a                                                                     : std_logic_vector(4 downto 0);   -- CPU_custom_instruction_master_multi_xconnect:ci_master0_a -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_n                                                                     : std_logic_vector(7 downto 0);   -- CPU_custom_instruction_master_multi_xconnect:ci_master0_n -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc                                                               : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_writerc -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending                                                              : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_xconnect:ci_master0_ipending -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk                                                                   : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_clk -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_start                                                                 : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_start -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa                                                                 : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_xconnect:ci_master0_dataa -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readra                                                                : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_readra -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_reset                                                                 : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_reset -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_datab                                                                 : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_xconnect:ci_master0_datab -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb                                                                : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_readrb -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus                                                               : std_logic;                      -- CPU_custom_instruction_master_multi_xconnect:ci_master0_estatus -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_result                                                        : std_logic_vector(31 downto 0);  -- nios_custom_instr_floating_point_0:result -> CPU_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_start                                                         : std_logic;                      -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_0:start
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa                                                         : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_0:dataa
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_done                                                          : std_logic;                      -- nios_custom_instr_floating_point_0:done -> CPU_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en                                                        : std_logic;                      -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_0:clk_en
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_n                                                             : std_logic_vector(1 downto 0);   -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_0:n
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset                                                         : std_logic;                      -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_0:reset
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab                                                         : std_logic_vector(31 downto 0);  -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_0:datab
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk                                                           : std_logic;                      -- CPU_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_0:clk
	signal cpu_instruction_master_waitrequest                                                                                            : std_logic;                      -- CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                                                                                : std_logic_vector(24 downto 0);  -- CPU:i_address -> CPU_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                                                   : std_logic;                      -- CPU:i_read -> CPU_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                                               : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	signal cpu_data_master_waitrequest                                                                                                   : std_logic;                      -- CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_writedata                                                                                                     : std_logic_vector(31 downto 0);  -- CPU:d_writedata -> CPU_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                                                       : std_logic_vector(24 downto 0);  -- CPU:d_address -> CPU_data_master_translator:av_address
	signal cpu_data_master_write                                                                                                         : std_logic;                      -- CPU:d_write -> CPU_data_master_translator:av_write
	signal cpu_data_master_read                                                                                                          : std_logic;                      -- CPU:d_read -> CPU_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                                                      : std_logic_vector(31 downto 0);  -- CPU_data_master_translator:av_readdata -> CPU:d_readdata
	signal cpu_data_master_debugaccess                                                                                                   : std_logic;                      -- CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                                                    : std_logic_vector(3 downto 0);   -- CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	signal pixel_buffer_dma_avalon_pixel_dma_master_waitrequest                                                                          : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_waitrequest -> Pixel_Buffer_DMA:master_waitrequest
	signal pixel_buffer_dma_avalon_pixel_dma_master_address                                                                              : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA:master_address -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_address
	signal pixel_buffer_dma_avalon_pixel_dma_master_lock                                                                                 : std_logic;                      -- Pixel_Buffer_DMA:master_arbiterlock -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_lock
	signal pixel_buffer_dma_avalon_pixel_dma_master_read                                                                                 : std_logic;                      -- Pixel_Buffer_DMA:master_read -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_read
	signal pixel_buffer_dma_avalon_pixel_dma_master_readdata                                                                             : std_logic_vector(7 downto 0);   -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_readdata -> Pixel_Buffer_DMA:master_readdata
	signal pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid                                                                        : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_readdatavalid -> Pixel_Buffer_DMA:master_readdatavalid
	signal video_dma_avalon_dma_master_waitrequest                                                                                       : std_logic;                      -- Video_DMA_avalon_dma_master_translator:av_waitrequest -> Video_DMA:master_waitrequest
	signal video_dma_avalon_dma_master_writedata                                                                                         : std_logic_vector(7 downto 0);   -- Video_DMA:master_writedata -> Video_DMA_avalon_dma_master_translator:av_writedata
	signal video_dma_avalon_dma_master_address                                                                                           : std_logic_vector(31 downto 0);  -- Video_DMA:master_address -> Video_DMA_avalon_dma_master_translator:av_address
	signal video_dma_avalon_dma_master_write                                                                                             : std_logic;                      -- Video_DMA:master_write -> Video_DMA_avalon_dma_master_translator:av_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                                              : std_logic;                      -- CPU:jtag_debug_module_waitrequest -> CPU_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                                                : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                                                  : std_logic_vector(8 downto 0);   -- CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                                                    : std_logic;                      -- CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                                                     : std_logic;                      -- CPU_jtag_debug_module_translator:av_read -> CPU:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                                              : std_logic;                      -- CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                                               : std_logic_vector(3 downto 0);   -- CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	signal onchip_memory_s1_translator_avalon_anti_slave_0_writedata                                                                     : std_logic_vector(31 downto 0);  -- Onchip_Memory_s1_translator:av_writedata -> Onchip_Memory:writedata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_address                                                                       : std_logic_vector(11 downto 0);  -- Onchip_Memory_s1_translator:av_address -> Onchip_Memory:address
	signal onchip_memory_s1_translator_avalon_anti_slave_0_chipselect                                                                    : std_logic;                      -- Onchip_Memory_s1_translator:av_chipselect -> Onchip_Memory:chipselect
	signal onchip_memory_s1_translator_avalon_anti_slave_0_clken                                                                         : std_logic;                      -- Onchip_Memory_s1_translator:av_clken -> Onchip_Memory:clken
	signal onchip_memory_s1_translator_avalon_anti_slave_0_write                                                                         : std_logic;                      -- Onchip_Memory_s1_translator:av_write -> Onchip_Memory:write
	signal onchip_memory_s1_translator_avalon_anti_slave_0_readdata                                                                      : std_logic_vector(31 downto 0);  -- Onchip_Memory:readdata -> Onchip_Memory_s1_translator:av_readdata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_byteenable                                                                    : std_logic_vector(3 downto 0);   -- Onchip_Memory_s1_translator:av_byteenable -> Onchip_Memory:byteenable
	signal sdram_0_s1_translator_avalon_anti_slave_0_waitrequest                                                                         : std_logic;                      -- sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	signal sdram_0_s1_translator_avalon_anti_slave_0_writedata                                                                           : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	signal sdram_0_s1_translator_avalon_anti_slave_0_address                                                                             : std_logic_vector(21 downto 0);  -- sdram_0_s1_translator:av_address -> sdram_0:az_addr
	signal sdram_0_s1_translator_avalon_anti_slave_0_chipselect                                                                          : std_logic;                      -- sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	signal sdram_0_s1_translator_avalon_anti_slave_0_write                                                                               : std_logic;                      -- sdram_0_s1_translator:av_write -> sdram_0_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_read                                                                                : std_logic;                      -- sdram_0_s1_translator:av_read -> sdram_0_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdata                                                                            : std_logic_vector(15 downto 0);  -- sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid                                                                       : std_logic;                      -- sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable                                                                          : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator:av_byteenable -> sdram_0_s1_translator_avalon_anti_slave_0_byteenable:in
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata                                                       : std_logic_vector(15 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator:av_writedata -> Pixel_Buffer:writedata
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address                                                         : std_logic_vector(17 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator:av_address -> Pixel_Buffer:address
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write                                                           : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator:av_write -> Pixel_Buffer:write
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read                                                            : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator:av_read -> Pixel_Buffer:read
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata                                                        : std_logic_vector(15 downto 0);  -- Pixel_Buffer:readdata -> Pixel_Buffer_avalon_sram_slave_translator:av_readdata
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid                                                   : std_logic;                      -- Pixel_Buffer:readdatavalid -> Pixel_Buffer_avalon_sram_slave_translator:av_readdatavalid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable                                                      : std_logic_vector(1 downto 0);   -- Pixel_Buffer_avalon_sram_slave_translator:av_byteenable -> Pixel_Buffer:byteenable
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest                                                   : std_logic;                      -- AV_Config:waitrequest -> AV_Config_avalon_av_config_slave_translator:av_waitrequest
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- AV_Config_avalon_av_config_slave_translator:av_writedata -> AV_Config:writedata
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- AV_Config_avalon_av_config_slave_translator:av_address -> AV_Config:address
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- AV_Config_avalon_av_config_slave_translator:av_write -> AV_Config:write
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read                                                          : std_logic;                      -- AV_Config_avalon_av_config_slave_translator:av_read -> AV_Config:read
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- AV_Config:readdata -> AV_Config_avalon_av_config_slave_translator:av_readdata
	signal av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable                                                    : std_logic_vector(3 downto 0);   -- AV_Config_avalon_av_config_slave_translator:av_byteenable -> AV_Config:byteenable
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- Video_DMA_avalon_dma_control_slave_translator:av_writedata -> Video_DMA:slave_writedata
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- Video_DMA_avalon_dma_control_slave_translator:av_address -> Video_DMA:slave_address
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator:av_write -> Video_DMA:slave_write
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read                                                        : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator:av_read -> Video_DMA:slave_read
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- Video_DMA:slave_readdata -> Video_DMA_avalon_dma_control_slave_translator:av_readdata
	signal video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable                                                  : std_logic_vector(3 downto 0);   -- Video_DMA_avalon_dma_control_slave_translator:av_byteenable -> Video_DMA:slave_byteenable
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA_avalon_control_slave_translator:av_writedata -> Pixel_Buffer_DMA:slave_writedata
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);   -- Pixel_Buffer_DMA_avalon_control_slave_translator:av_address -> Pixel_Buffer_DMA:slave_address
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write                                                    : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator:av_write -> Pixel_Buffer_DMA:slave_write
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read                                                     : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator:av_read -> Pixel_Buffer_DMA:slave_read
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA:slave_readdata -> Pixel_Buffer_DMA_avalon_control_slave_translator:av_readdata
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable                                               : std_logic_vector(3 downto 0);   -- Pixel_Buffer_DMA_avalon_control_slave_translator:av_byteenable -> Pixel_Buffer_DMA:slave_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                                      : std_logic;                      -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                                        : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                                          : std_logic_vector(0 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                                            : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                                             : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                                         : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address                                                             : std_logic_vector(0 downto 0);   -- sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata                                                            : std_logic_vector(31 downto 0);  -- sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	signal timer_system_s1_translator_avalon_anti_slave_0_writedata                                                                      : std_logic_vector(15 downto 0);  -- timer_system_s1_translator:av_writedata -> timer_system:writedata
	signal timer_system_s1_translator_avalon_anti_slave_0_address                                                                        : std_logic_vector(2 downto 0);   -- timer_system_s1_translator:av_address -> timer_system:address
	signal timer_system_s1_translator_avalon_anti_slave_0_chipselect                                                                     : std_logic;                      -- timer_system_s1_translator:av_chipselect -> timer_system:chipselect
	signal timer_system_s1_translator_avalon_anti_slave_0_write                                                                          : std_logic;                      -- timer_system_s1_translator:av_write -> timer_system_s1_translator_avalon_anti_slave_0_write:in
	signal timer_system_s1_translator_avalon_anti_slave_0_readdata                                                                       : std_logic_vector(15 downto 0);  -- timer_system:readdata -> timer_system_s1_translator:av_readdata
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_writedata                                                                   : std_logic_vector(15 downto 0);  -- timer_timestamp_s1_translator:av_writedata -> timer_timestamp:writedata
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_address                                                                     : std_logic_vector(2 downto 0);   -- timer_timestamp_s1_translator:av_address -> timer_timestamp:address
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect                                                                  : std_logic;                      -- timer_timestamp_s1_translator:av_chipselect -> timer_timestamp:chipselect
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_write                                                                       : std_logic;                      -- timer_timestamp_s1_translator:av_write -> timer_timestamp_s1_translator_avalon_anti_slave_0_write:in
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_readdata                                                                    : std_logic_vector(15 downto 0);  -- timer_timestamp:readdata -> timer_timestamp_s1_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_writedata                                                                    : std_logic_vector(7 downto 0);   -- lcd_control_slave_translator:av_writedata -> lcd:writedata
	signal lcd_control_slave_translator_avalon_anti_slave_0_address                                                                      : std_logic_vector(1 downto 0);   -- lcd_control_slave_translator:av_address -> lcd:address
	signal lcd_control_slave_translator_avalon_anti_slave_0_write                                                                        : std_logic;                      -- lcd_control_slave_translator:av_write -> lcd:write
	signal lcd_control_slave_translator_avalon_anti_slave_0_read                                                                         : std_logic;                      -- lcd_control_slave_translator:av_read -> lcd:read
	signal lcd_control_slave_translator_avalon_anti_slave_0_readdata                                                                     : std_logic_vector(7 downto 0);   -- lcd:readdata -> lcd_control_slave_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_begintransfer                                                                : std_logic;                      -- lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	signal red_leds_s1_translator_avalon_anti_slave_0_writedata                                                                          : std_logic_vector(31 downto 0);  -- red_leds_s1_translator:av_writedata -> red_leds:writedata
	signal red_leds_s1_translator_avalon_anti_slave_0_address                                                                            : std_logic_vector(1 downto 0);   -- red_leds_s1_translator:av_address -> red_leds:address
	signal red_leds_s1_translator_avalon_anti_slave_0_chipselect                                                                         : std_logic;                      -- red_leds_s1_translator:av_chipselect -> red_leds:chipselect
	signal red_leds_s1_translator_avalon_anti_slave_0_write                                                                              : std_logic;                      -- red_leds_s1_translator:av_write -> red_leds_s1_translator_avalon_anti_slave_0_write:in
	signal red_leds_s1_translator_avalon_anti_slave_0_readdata                                                                           : std_logic_vector(31 downto 0);  -- red_leds:readdata -> red_leds_s1_translator:av_readdata
	signal green_leds_s1_translator_avalon_anti_slave_0_writedata                                                                        : std_logic_vector(31 downto 0);  -- green_leds_s1_translator:av_writedata -> green_leds:writedata
	signal green_leds_s1_translator_avalon_anti_slave_0_address                                                                          : std_logic_vector(1 downto 0);   -- green_leds_s1_translator:av_address -> green_leds:address
	signal green_leds_s1_translator_avalon_anti_slave_0_chipselect                                                                       : std_logic;                      -- green_leds_s1_translator:av_chipselect -> green_leds:chipselect
	signal green_leds_s1_translator_avalon_anti_slave_0_write                                                                            : std_logic;                      -- green_leds_s1_translator:av_write -> green_leds_s1_translator_avalon_anti_slave_0_write:in
	signal green_leds_s1_translator_avalon_anti_slave_0_readdata                                                                         : std_logic_vector(31 downto 0);  -- green_leds:readdata -> green_leds_s1_translator:av_readdata
	signal switch_s1_translator_avalon_anti_slave_0_address                                                                              : std_logic_vector(1 downto 0);   -- switch_s1_translator:av_address -> switch:address
	signal switch_s1_translator_avalon_anti_slave_0_readdata                                                                             : std_logic_vector(31 downto 0);  -- switch:readdata -> switch_s1_translator:av_readdata
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_waitrequest
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(7 downto 0);   -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_readdata
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_writedata                                                                    : std_logic_vector(7 downto 0);   -- Barcode_scan_0_s1_translator:av_writedata -> Barcode_scan_0:avs_s1_writedata
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_address                                                                      : std_logic_vector(7 downto 0);   -- Barcode_scan_0_s1_translator:av_address -> Barcode_scan_0:avs_s1_address
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_chipselect                                                                   : std_logic;                      -- Barcode_scan_0_s1_translator:av_chipselect -> Barcode_scan_0:avs_s1_chipselect
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_write                                                                        : std_logic;                      -- Barcode_scan_0_s1_translator:av_write -> Barcode_scan_0:avs_s1_write
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_read                                                                         : std_logic;                      -- Barcode_scan_0_s1_translator:av_read -> Barcode_scan_0:avs_s1_read
	signal barcode_scan_0_s1_translator_avalon_anti_slave_0_readdata                                                                     : std_logic_vector(7 downto 0);   -- Barcode_scan_0:avs_s1_readdata -> Barcode_scan_0_s1_translator:av_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                                                       : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                                                        : std_logic_vector(2 downto 0);   -- CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                                                         : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                                                           : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                                              : std_logic;                      -- CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                                             : std_logic;                      -- CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                                              : std_logic;                      -- CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                                                          : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                                                       : std_logic;                      -- CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                                                        : std_logic_vector(3 downto 0);   -- CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                                                     : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                                              : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                                               : std_logic_vector(2 downto 0);   -- CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                                                : std_logic_vector(31 downto 0);  -- CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                                                  : std_logic_vector(31 downto 0);  -- CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                                                     : std_logic;                      -- CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                                                    : std_logic;                      -- CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                                                     : std_logic;                      -- CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                                                 : std_logic_vector(31 downto 0);  -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                                              : std_logic;                      -- CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                                               : std_logic_vector(3 downto 0);   -- CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                                                            : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest                                     : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_waitrequest
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount                                      : std_logic_vector(0 downto 0);   -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_burstcount -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata                                       : std_logic_vector(7 downto 0);   -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_writedata -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address                                         : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_address -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock                                            : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_lock -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write                                           : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_write -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read                                            : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_read -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata                                        : std_logic_vector(7 downto 0);   -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_readdata
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess                                     : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_debugaccess -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable                                      : std_logic_vector(0 downto 0);   -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_byteenable -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid                                   : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_readdatavalid
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest                                                  : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Video_DMA_avalon_dma_master_translator:uav_waitrequest
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount                                                   : std_logic_vector(0 downto 0);   -- Video_DMA_avalon_dma_master_translator:uav_burstcount -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata                                                    : std_logic_vector(7 downto 0);   -- Video_DMA_avalon_dma_master_translator:uav_writedata -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_address                                                      : std_logic_vector(31 downto 0);  -- Video_DMA_avalon_dma_master_translator:uav_address -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock                                                         : std_logic;                      -- Video_DMA_avalon_dma_master_translator:uav_lock -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_write                                                        : std_logic;                      -- Video_DMA_avalon_dma_master_translator:uav_write -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_read                                                         : std_logic;                      -- Video_DMA_avalon_dma_master_translator:uav_read -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata                                                     : std_logic_vector(7 downto 0);   -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Video_DMA_avalon_dma_master_translator:uav_readdata
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess                                                  : std_logic;                      -- Video_DMA_avalon_dma_master_translator:uav_debugaccess -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable                                                   : std_logic_vector(0 downto 0);   -- Video_DMA_avalon_dma_master_translator:uav_byteenable -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid                                                : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Video_DMA_avalon_dma_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                : std_logic;                      -- CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                                                 : std_logic_vector(2 downto 0);   -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                                                  : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                                                    : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                                                      : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                                                       : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                                                       : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                                                   : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                              : std_logic;                      -- CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                                                 : std_logic_vector(3 downto 0);   -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                         : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                                               : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                       : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                                                : std_logic_vector(109 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                                               : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                      : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                            : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                    : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                             : std_logic_vector(109 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                            : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                          : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                           : std_logic_vector(33 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                          : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                     : std_logic;                      -- Onchip_Memory_s1_translator:uav_waitrequest -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                      : std_logic_vector(2 downto 0);   -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_Memory_s1_translator:uav_burstcount
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                       : std_logic_vector(31 downto 0);  -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_Memory_s1_translator:uav_writedata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                                                         : std_logic_vector(31 downto 0);  -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_Memory_s1_translator:uav_address
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                                                           : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_Memory_s1_translator:uav_write
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                            : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_Memory_s1_translator:uav_lock
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                                            : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_Memory_s1_translator:uav_read
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                        : std_logic_vector(31 downto 0);  -- Onchip_Memory_s1_translator:uav_readdata -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                   : std_logic;                      -- Onchip_Memory_s1_translator:uav_readdatavalid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                     : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_Memory_s1_translator:uav_debugaccess
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                      : std_logic_vector(3 downto 0);   -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_Memory_s1_translator:uav_byteenable
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                              : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                    : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                            : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                     : std_logic_vector(109 downto 0); -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                    : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                           : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                 : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                         : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                  : std_logic_vector(109 downto 0); -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                 : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                               : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                : std_logic_vector(33 downto 0);  -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                               : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                           : std_logic;                      -- sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                            : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                             : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                               : std_logic_vector(31 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                                 : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                              : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                         : std_logic;                      -- sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                            : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                                    : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                           : std_logic_vector(91 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                                 : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                       : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                               : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                        : std_logic_vector(91 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                       : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                                     : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                      : std_logic_vector(17 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                                     : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                                     : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                                      : std_logic_vector(17 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                                     : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                       : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator:uav_waitrequest -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                        : std_logic_vector(1 downto 0);   -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pixel_Buffer_avalon_sram_slave_translator:uav_burstcount
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                         : std_logic_vector(15 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pixel_Buffer_avalon_sram_slave_translator:uav_writedata
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address                                           : std_logic_vector(31 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pixel_Buffer_avalon_sram_slave_translator:uav_address
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write                                             : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pixel_Buffer_avalon_sram_slave_translator:uav_write
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock                                              : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pixel_Buffer_avalon_sram_slave_translator:uav_lock
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read                                              : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pixel_Buffer_avalon_sram_slave_translator:uav_read
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                          : std_logic_vector(15 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator:uav_readdata -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                     : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator:uav_readdatavalid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                       : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pixel_Buffer_avalon_sram_slave_translator:uav_debugaccess
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                        : std_logic_vector(1 downto 0);   -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pixel_Buffer_avalon_sram_slave_translator:uav_byteenable
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                      : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                              : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                       : std_logic_vector(91 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                      : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                             : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                   : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                           : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                    : std_logic_vector(91 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                   : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                 : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                  : std_logic_vector(17 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                 : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                 : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                  : std_logic_vector(17 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                 : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- AV_Config_avalon_av_config_slave_translator:uav_waitrequest -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> AV_Config_avalon_av_config_slave_translator:uav_burstcount
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> AV_Config_avalon_av_config_slave_translator:uav_writedata
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(31 downto 0);  -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> AV_Config_avalon_av_config_slave_translator:uav_address
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> AV_Config_avalon_av_config_slave_translator:uav_write
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> AV_Config_avalon_av_config_slave_translator:uav_lock
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> AV_Config_avalon_av_config_slave_translator:uav_read
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- AV_Config_avalon_av_config_slave_translator:uav_readdata -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- AV_Config_avalon_av_config_slave_translator:uav_readdatavalid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> AV_Config_avalon_av_config_slave_translator:uav_debugaccess
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> AV_Config_avalon_av_config_slave_translator:uav_byteenable
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(109 downto 0); -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(109 downto 0); -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator:uav_waitrequest -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Video_DMA_avalon_dma_control_slave_translator:uav_burstcount
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Video_DMA_avalon_dma_control_slave_translator:uav_writedata
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(31 downto 0);  -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Video_DMA_avalon_dma_control_slave_translator:uav_address
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Video_DMA_avalon_dma_control_slave_translator:uav_write
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Video_DMA_avalon_dma_control_slave_translator:uav_lock
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Video_DMA_avalon_dma_control_slave_translator:uav_read
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- Video_DMA_avalon_dma_control_slave_translator:uav_readdata -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator:uav_readdatavalid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Video_DMA_avalon_dma_control_slave_translator:uav_debugaccess
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Video_DMA_avalon_dma_control_slave_translator:uav_byteenable
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(109 downto 0); -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(109 downto 0); -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator:uav_waitrequest -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);   -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_burstcount
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_writedata
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_address
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_write
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_lock
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_read
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0);  -- Pixel_Buffer_DMA_avalon_control_slave_translator:uav_readdata -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator:uav_readdatavalid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_debugaccess
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);   -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_byteenable
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(109 downto 0); -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(109 downto 0); -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0);  -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                         : std_logic_vector(2 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                          : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                                            : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                           : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                         : std_logic_vector(3 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                        : std_logic_vector(109 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                    : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                            : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                     : std_logic_vector(109 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                    : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                   : std_logic_vector(33 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                           : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                            : std_logic_vector(2 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                             : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                               : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                              : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                         : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                            : std_logic_vector(3 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                    : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                          : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                           : std_logic_vector(109 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                          : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                       : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                               : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                        : std_logic_vector(109 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                       : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                     : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                      : std_logic_vector(33 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                     : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                      : std_logic;                      -- timer_system_s1_translator:uav_waitrequest -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                       : std_logic_vector(2 downto 0);   -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_system_s1_translator:uav_burstcount
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                        : std_logic_vector(31 downto 0);  -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_system_s1_translator:uav_writedata
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address                                                          : std_logic_vector(31 downto 0);  -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_system_s1_translator:uav_address
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write                                                            : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_system_s1_translator:uav_write
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                             : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_system_s1_translator:uav_lock
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read                                                             : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_system_s1_translator:uav_read
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                         : std_logic_vector(31 downto 0);  -- timer_system_s1_translator:uav_readdata -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                    : std_logic;                      -- timer_system_s1_translator:uav_readdatavalid -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                      : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_system_s1_translator:uav_debugaccess
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                       : std_logic_vector(3 downto 0);   -- timer_system_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_system_s1_translator:uav_byteenable
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                               : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                     : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                             : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                      : std_logic_vector(109 downto 0); -- timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                     : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                            : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                  : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                          : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                   : std_logic_vector(109 downto 0); -- timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                  : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                                : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                 : std_logic_vector(33 downto 0);  -- timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                                : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                   : std_logic;                      -- timer_timestamp_s1_translator:uav_waitrequest -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                    : std_logic_vector(2 downto 0);   -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_timestamp_s1_translator:uav_burstcount
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                     : std_logic_vector(31 downto 0);  -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_timestamp_s1_translator:uav_writedata
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address                                                       : std_logic_vector(31 downto 0);  -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_timestamp_s1_translator:uav_address
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write                                                         : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_timestamp_s1_translator:uav_write
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                          : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_timestamp_s1_translator:uav_lock
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read                                                          : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_timestamp_s1_translator:uav_read
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                      : std_logic_vector(31 downto 0);  -- timer_timestamp_s1_translator:uav_readdata -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                 : std_logic;                      -- timer_timestamp_s1_translator:uav_readdatavalid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                   : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_timestamp_s1_translator:uav_debugaccess
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                    : std_logic_vector(3 downto 0);   -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_timestamp_s1_translator:uav_byteenable
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                            : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                  : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                          : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                   : std_logic_vector(109 downto 0); -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                  : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                         : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                               : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                       : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                : std_logic_vector(109 downto 0); -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                               : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                             : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                              : std_logic_vector(33 downto 0);  -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                             : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                    : std_logic;                      -- lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                                     : std_logic_vector(2 downto 0);   -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                                      : std_logic_vector(31 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                                        : std_logic_vector(31 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                                          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                                           : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                                           : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                                       : std_logic_vector(31 downto 0);  -- lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                  : std_logic;                      -- lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                    : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                                     : std_logic_vector(3 downto 0);   -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                             : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                                                   : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                           : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                                                    : std_logic_vector(109 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                                                   : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                        : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                 : std_logic_vector(109 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                              : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                               : std_logic_vector(33 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                              : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                          : std_logic;                      -- red_leds_s1_translator:uav_waitrequest -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                           : std_logic_vector(2 downto 0);   -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> red_leds_s1_translator:uav_burstcount
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                            : std_logic_vector(31 downto 0);  -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> red_leds_s1_translator:uav_writedata
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address                                                              : std_logic_vector(31 downto 0);  -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> red_leds_s1_translator:uav_address
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write                                                                : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> red_leds_s1_translator:uav_write
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                                 : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> red_leds_s1_translator:uav_lock
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read                                                                 : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> red_leds_s1_translator:uav_read
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                             : std_logic_vector(31 downto 0);  -- red_leds_s1_translator:uav_readdata -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                        : std_logic;                      -- red_leds_s1_translator:uav_readdatavalid -> red_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                          : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> red_leds_s1_translator:uav_debugaccess
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                           : std_logic_vector(3 downto 0);   -- red_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> red_leds_s1_translator:uav_byteenable
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                                   : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                         : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                                 : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                          : std_logic_vector(109 downto 0); -- red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                         : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                                : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                      : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                              : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                       : std_logic_vector(109 downto 0); -- red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                      : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                                    : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                     : std_logic_vector(33 downto 0);  -- red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                                    : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                        : std_logic;                      -- green_leds_s1_translator:uav_waitrequest -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                         : std_logic_vector(2 downto 0);   -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_leds_s1_translator:uav_burstcount
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                          : std_logic_vector(31 downto 0);  -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_leds_s1_translator:uav_writedata
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address                                                            : std_logic_vector(31 downto 0);  -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_leds_s1_translator:uav_address
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write                                                              : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_leds_s1_translator:uav_write
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                               : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_leds_s1_translator:uav_lock
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read                                                               : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_leds_s1_translator:uav_read
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                           : std_logic_vector(31 downto 0);  -- green_leds_s1_translator:uav_readdata -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                      : std_logic;                      -- green_leds_s1_translator:uav_readdatavalid -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                        : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_leds_s1_translator:uav_debugaccess
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                         : std_logic_vector(3 downto 0);   -- green_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_leds_s1_translator:uav_byteenable
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                                 : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                       : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                               : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                        : std_logic_vector(109 downto 0); -- green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                       : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                              : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                    : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                            : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                     : std_logic_vector(109 downto 0); -- green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                    : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                                  : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                   : std_logic_vector(33 downto 0);  -- green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                                  : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                            : std_logic;                      -- switch_s1_translator:uav_waitrequest -> switch_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                             : std_logic_vector(2 downto 0);   -- switch_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_s1_translator:uav_burstcount
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                              : std_logic_vector(31 downto 0);  -- switch_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_s1_translator:uav_writedata
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_address                                                                : std_logic_vector(31 downto 0);  -- switch_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_s1_translator:uav_address
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_write                                                                  : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_s1_translator:uav_write
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                                   : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_s1_translator:uav_lock
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_read                                                                   : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_s1_translator:uav_read
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                               : std_logic_vector(31 downto 0);  -- switch_s1_translator:uav_readdata -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                          : std_logic;                      -- switch_s1_translator:uav_readdatavalid -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                            : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_s1_translator:uav_debugaccess
	signal switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                             : std_logic_vector(3 downto 0);   -- switch_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_s1_translator:uav_byteenable
	signal switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                                     : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                           : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                                   : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                            : std_logic_vector(109 downto 0); -- switch_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                           : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                                  : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                        : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                                : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                         : std_logic_vector(109 downto 0); -- switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                        : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                                      : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                                       : std_logic_vector(33 downto 0);  -- switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                                      : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_burstcount
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_writedata
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_address
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_write
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_lock
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_read
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdatavalid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_debugaccess
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_byteenable
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(109 downto 0); -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(109 downto 0); -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                                    : std_logic;                      -- Barcode_scan_0_s1_translator:uav_waitrequest -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                                     : std_logic_vector(0 downto 0);   -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Barcode_scan_0_s1_translator:uav_burstcount
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                                      : std_logic_vector(7 downto 0);   -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Barcode_scan_0_s1_translator:uav_writedata
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                                        : std_logic_vector(31 downto 0);  -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> Barcode_scan_0_s1_translator:uav_address
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                                          : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> Barcode_scan_0_s1_translator:uav_write
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                           : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Barcode_scan_0_s1_translator:uav_lock
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                                           : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> Barcode_scan_0_s1_translator:uav_read
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                                       : std_logic_vector(7 downto 0);   -- Barcode_scan_0_s1_translator:uav_readdata -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                                  : std_logic;                      -- Barcode_scan_0_s1_translator:uav_readdatavalid -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                                    : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Barcode_scan_0_s1_translator:uav_debugaccess
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                                     : std_logic_vector(0 downto 0);   -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Barcode_scan_0_s1_translator:uav_byteenable
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                             : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                                   : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                           : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                                    : std_logic_vector(82 downto 0);  -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                                   : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                          : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                                : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                        : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                                 : std_logic_vector(82 downto 0);  -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                                : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                              : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                               : std_logic_vector(9 downto 0);   -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                              : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                              : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                                                    : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                            : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                                                     : std_logic_vector(108 downto 0); -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                                                    : std_logic;                      -- addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                                     : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                                                           : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                                   : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                                                            : std_logic_vector(108 downto 0); -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                                                           : std_logic;                      -- addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket                            : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid                                  : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket                          : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data                                   : std_logic_vector(81 downto 0);  -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready                                  : std_logic;                      -- addr_router_002:sink_ready -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                         : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid                                               : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                       : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data                                                : std_logic_vector(81 downto 0);  -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	signal video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready                                               : std_logic;                      -- addr_router_003:sink_ready -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                                                      : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                                              : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                                                       : std_logic_vector(108 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                                                      : std_logic;                      -- id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                     : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                           : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                   : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                                            : std_logic_vector(108 downto 0); -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                           : std_logic;                      -- id_router_001:sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                                 : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                         : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                                  : std_logic_vector(90 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                                 : std_logic;                      -- id_router_002:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                       : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid                                             : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                     : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data                                              : std_logic_vector(90 downto 0);  -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready                                             : std_logic;                      -- id_router_003:sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(108 downto 0); -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_004:sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(108 downto 0); -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_005:sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(108 downto 0); -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                      -- id_router_006:sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                                              : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                                               : std_logic_vector(108 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                                              : std_logic;                      -- id_router_007:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                         : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                                  : std_logic_vector(108 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                                 : std_logic;                      -- id_router_008:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                      : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                            : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                    : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data                                                             : std_logic_vector(108 downto 0); -- timer_system_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                            : std_logic;                      -- id_router_009:sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                   : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                         : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                 : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data                                                          : std_logic_vector(108 downto 0); -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                         : std_logic;                      -- id_router_010:sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                    : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                                          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                  : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                                           : std_logic_vector(108 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                                          : std_logic;                      -- id_router_011:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                          : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                                : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                        : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data                                                                 : std_logic_vector(108 downto 0); -- red_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                                : std_logic;                      -- id_router_012:sink_ready -> red_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                        : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                              : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                      : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data                                                               : std_logic_vector(108 downto 0); -- green_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                              : std_logic;                      -- id_router_013:sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                            : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                                  : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                          : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal switch_s1_translator_avalon_universal_slave_0_agent_rp_data                                                                   : std_logic_vector(108 downto 0); -- switch_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal switch_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                                  : std_logic;                      -- id_router_014:sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(108 downto 0); -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_015:sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                                    : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                          : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                                  : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                                           : std_logic_vector(81 downto 0);  -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                          : std_logic;                      -- id_router_016:sink_ready -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                                                             : std_logic;                      -- burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                                                   : std_logic;                      -- burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                                           : std_logic;                      -- burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                                                    : std_logic_vector(90 downto 0);  -- burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                                                   : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                                                 : std_logic_vector(16 downto 0);  -- burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                                         : std_logic;                      -- burst_adapter_001:source0_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                                               : std_logic;                      -- burst_adapter_001:source0_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                                                       : std_logic;                      -- burst_adapter_001:source0_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                                                : std_logic_vector(90 downto 0);  -- burst_adapter_001:source0_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                                               : std_logic;                      -- Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                                             : std_logic_vector(16 downto 0);  -- burst_adapter_001:source0_channel -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_002_source0_endofpacket                                                                                         : std_logic;                      -- burst_adapter_002:source0_endofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_002_source0_valid                                                                                               : std_logic;                      -- burst_adapter_002:source0_valid -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_002_source0_startofpacket                                                                                       : std_logic;                      -- burst_adapter_002:source0_startofpacket -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_002_source0_data                                                                                                : std_logic_vector(81 downto 0);  -- burst_adapter_002:source0_data -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_002_source0_ready                                                                                               : std_logic;                      -- Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	signal burst_adapter_002_source0_channel                                                                                             : std_logic_vector(16 downto 0);  -- burst_adapter_002:source0_channel -> Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                                                : std_logic;                      -- rst_controller:reset_out -> [AV_Config:reset, AV_Config_avalon_av_config_slave_translator:reset, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Barcode_scan_0_s1_translator:reset, Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent:reset, Barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Dual_Clock_FIFO:reset_stream_in, Onchip_Memory:reset, Onchip_Memory_s1_translator:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_Buffer:reset, Pixel_Buffer_DMA:reset, Pixel_Buffer_DMA_avalon_control_slave_translator:reset, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:reset, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, Pixel_Buffer_avalon_sram_slave_translator:reset, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_RGB_Resampler:reset, Video_DMA:reset, Video_DMA_avalon_dma_control_slave_translator:reset, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Video_DMA_avalon_dma_master_translator:reset, Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, Video_In_Decoder:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, green_leds_s1_translator:reset, green_leds_s1_translator_avalon_universal_slave_0_agent:reset, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, red_leds_s1_translator:reset, red_leds_s1_translator_avalon_universal_slave_0_agent:reset, red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch_s1_translator:reset, switch_s1_translator_avalon_universal_slave_0_agent:reset, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_system_s1_translator:reset, timer_system_s1_translator_avalon_universal_slave_0_agent:reset, timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_timestamp_s1_translator:reset, timer_timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_bayer_resampler:reset, video_clipper_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset]
	signal rst_controller_reset_out_reset_req                                                                                            : std_logic;                      -- rst_controller:reset_req -> Onchip_Memory:reset_req
	signal cpu_jtag_debug_module_reset_reset                                                                                             : std_logic;                      -- CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal clock_signals_sys_clk_reset_reset                                                                                             : std_logic;                      -- Clock_Signals:sys_reset_n -> clock_signals_sys_clk_reset_reset:in
	signal rst_controller_001_reset_out_reset                                                                                            : std_logic;                      -- rst_controller_001:reset_out -> [Dual_Clock_FIFO:reset_stream_out, VGA_Controller:reset]
	signal rst_controller_002_reset_out_reset                                                                                            : std_logic;                      -- rst_controller_002:reset_out -> Clock_Signals:reset
	signal rst_controller_003_reset_out_reset                                                                                            : std_logic;                      -- rst_controller_003:reset_out -> [rst_controller:reset_in3, rst_controller_001:reset_in3, rst_controller_002:reset_in3]
	signal cmd_xbar_demux_src0_endofpacket                                                                                               : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                                     : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                                             : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                                      : std_logic_vector(108 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                                                   : std_logic_vector(16 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                                     : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                                               : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                                     : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                                             : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                                      : std_logic_vector(108 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                                                   : std_logic_vector(16 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                                                     : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                                                 : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                                                 : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src4_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src4_channel -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src5_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src5_channel -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src6_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src6_channel -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src7_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src7_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src8_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src8_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src9_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src9_channel -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src10_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src10_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src10_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src10_channel -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src11_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src11_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src11_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src11_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src11_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src11_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src11_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src12_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src12_endofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src12_valid -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src12_startofpacket -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src12_data -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src12_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src12_channel -> red_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src13_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src13_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src13_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src13_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src13_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src13_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src13_channel -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src14_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src14_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src14_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src14_valid -> switch_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src14_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src14_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src14_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src14_data -> switch_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src14_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src14_channel -> switch_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src15_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src15_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src15_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src15_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src15_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src15_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src15_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src15_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src15_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src15_channel -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                                               : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                                     : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                                             : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                                      : std_logic_vector(108 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                                                   : std_logic_vector(16 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                                     : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                                               : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                                     : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                                             : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                                      : std_logic_vector(108 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                                                   : std_logic_vector(16 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                                     : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                                                  : std_logic_vector(108 downto 0); -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	signal rsp_xbar_demux_015_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	signal rsp_xbar_demux_015_src0_ready                                                                                                 : std_logic;                      -- rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	signal addr_router_src_endofpacket                                                                                                   : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                                         : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                                                 : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                                          : std_logic_vector(108 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                                       : std_logic_vector(16 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                                         : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                                                  : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                                        : std_logic;                      -- rsp_xbar_mux:src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                                                : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                                         : std_logic_vector(108 downto 0); -- rsp_xbar_mux:src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                                                      : std_logic_vector(16 downto 0);  -- rsp_xbar_mux:src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                                        : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                                               : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                                     : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                                             : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                                      : std_logic_vector(108 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                                                   : std_logic_vector(16 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                                     : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                                              : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                                                    : std_logic;                      -- rsp_xbar_mux_001:src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                                            : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                                                     : std_logic_vector(108 downto 0); -- rsp_xbar_mux_001:src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                                                  : std_logic_vector(16 downto 0);  -- rsp_xbar_mux_001:src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                                                    : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal addr_router_002_src_endofpacket                                                                                               : std_logic;                      -- addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal addr_router_002_src_valid                                                                                                     : std_logic;                      -- addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	signal addr_router_002_src_startofpacket                                                                                             : std_logic;                      -- addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal addr_router_002_src_data                                                                                                      : std_logic_vector(81 downto 0);  -- addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	signal addr_router_002_src_channel                                                                                                   : std_logic_vector(16 downto 0);  -- addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	signal addr_router_002_src_ready                                                                                                     : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	signal width_adapter_009_src_ready                                                                                                   : std_logic;                      -- Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_009:out_ready
	signal addr_router_003_src_endofpacket                                                                                               : std_logic;                      -- addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	signal addr_router_003_src_valid                                                                                                     : std_logic;                      -- addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	signal addr_router_003_src_startofpacket                                                                                             : std_logic;                      -- addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	signal addr_router_003_src_data                                                                                                      : std_logic_vector(81 downto 0);  -- addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	signal addr_router_003_src_channel                                                                                                   : std_logic_vector(16 downto 0);  -- addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	signal addr_router_003_src_ready                                                                                                     : std_logic;                      -- cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	signal width_adapter_010_src_ready                                                                                                   : std_logic;                      -- Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_010:out_ready
	signal cmd_xbar_mux_src_endofpacket                                                                                                  : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                                        : std_logic;                      -- cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                                                : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                                         : std_logic_vector(108 downto 0); -- cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                                      : std_logic_vector(16 downto 0);  -- cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                                        : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                                     : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                                           : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                                                   : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                                            : std_logic_vector(108 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                                         : std_logic_vector(16 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                                           : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                                              : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                                                    : std_logic;                      -- cmd_xbar_mux_001:src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                                            : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                                                     : std_logic_vector(108 downto 0); -- cmd_xbar_mux_001:src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                                                  : std_logic_vector(16 downto 0);  -- cmd_xbar_mux_001:src_channel -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                                                    : std_logic;                      -- Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                                                 : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                                       : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                                               : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                                              : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                                                    : std_logic;                      -- cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                                            : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                                                     : std_logic_vector(90 downto 0);  -- cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_002_src_channel                                                                                                  : std_logic_vector(16 downto 0);  -- cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_002_src_ready                                                                                                    : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                                                 : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                                       : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                                               : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                                        : std_logic_vector(90 downto 0);  -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                                              : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                                                    : std_logic;                      -- cmd_xbar_mux_003:src_valid -> burst_adapter_001:sink0_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                                            : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                                                     : std_logic_vector(90 downto 0);  -- cmd_xbar_mux_003:src_data -> burst_adapter_001:sink0_data
	signal cmd_xbar_mux_003_src_channel                                                                                                  : std_logic_vector(16 downto 0);  -- cmd_xbar_mux_003:src_channel -> burst_adapter_001:sink0_channel
	signal cmd_xbar_mux_003_src_ready                                                                                                    : std_logic;                      -- burst_adapter_001:sink0_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                                                 : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                                       : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                                               : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                                        : std_logic_vector(90 downto 0);  -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                                                 : std_logic;                      -- AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                                                 : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                                       : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                                               : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                                                 : std_logic;                      -- Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                                                 : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                                       : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                                               : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                                                 : std_logic;                      -- Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                                                 : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                                       : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                                               : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                                                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                                                 : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                                       : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                                               : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                                                 : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                                                 : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                                       : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                                               : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                                                 : std_logic;                      -- timer_system_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                                                 : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                                       : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                                               : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_001_src10_ready                                                                                                : std_logic;                      -- timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	signal id_router_010_src_endofpacket                                                                                                 : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                                       : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                                               : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_001_src11_ready                                                                                                : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	signal id_router_011_src_endofpacket                                                                                                 : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                                                       : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                                               : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_001_src12_ready                                                                                                : std_logic;                      -- red_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	signal id_router_012_src_endofpacket                                                                                                 : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                                                       : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                                               : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_001_src13_ready                                                                                                : std_logic;                      -- green_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	signal id_router_013_src_endofpacket                                                                                                 : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                                                       : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                                               : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_demux_001_src14_ready                                                                                                : std_logic;                      -- switch_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	signal id_router_014_src_endofpacket                                                                                                 : std_logic;                      -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                                                       : std_logic;                      -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                                                               : std_logic;                      -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_demux_001_src15_ready                                                                                                : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	signal id_router_015_src_endofpacket                                                                                                 : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                                                       : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                                               : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                                                        : std_logic_vector(108 downto 0); -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal width_adapter_003_src_ready                                                                                                   : std_logic;                      -- burst_adapter_002:sink0_ready -> width_adapter_003:out_ready
	signal id_router_016_src_endofpacket                                                                                                 : std_logic;                      -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                                                       : std_logic;                      -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                                                               : std_logic;                      -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                                                        : std_logic_vector(81 downto 0);  -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                                                       : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                                               : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                                                     : std_logic;                      -- cmd_xbar_demux:src2_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                                             : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src2_data                                                                                                      : std_logic_vector(108 downto 0); -- cmd_xbar_demux:src2_data -> width_adapter:in_data
	signal cmd_xbar_demux_src2_channel                                                                                                   : std_logic_vector(16 downto 0);  -- cmd_xbar_demux:src2_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_src2_ready                                                                                                     : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux:src2_ready
	signal width_adapter_src_endofpacket                                                                                                 : std_logic;                      -- width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal width_adapter_src_valid                                                                                                       : std_logic;                      -- width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	signal width_adapter_src_startofpacket                                                                                               : std_logic;                      -- width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal width_adapter_src_data                                                                                                        : std_logic_vector(90 downto 0);  -- width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	signal width_adapter_src_ready                                                                                                       : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                                                     : std_logic_vector(16 downto 0);  -- width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_001_src2_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> width_adapter_001:in_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> width_adapter_001:in_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> width_adapter_001:in_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src2_data -> width_adapter_001:in_data
	signal cmd_xbar_demux_001_src2_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src2_channel -> width_adapter_001:in_channel
	signal cmd_xbar_demux_001_src2_ready                                                                                                 : std_logic;                      -- width_adapter_001:in_ready -> cmd_xbar_demux_001:src2_ready
	signal width_adapter_001_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal width_adapter_001_src_valid                                                                                                   : std_logic;                      -- width_adapter_001:out_valid -> cmd_xbar_mux_002:sink1_valid
	signal width_adapter_001_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal width_adapter_001_src_data                                                                                                    : std_logic_vector(90 downto 0);  -- width_adapter_001:out_data -> cmd_xbar_mux_002:sink1_data
	signal width_adapter_001_src_ready                                                                                                   : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_001:out_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                                                  : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src3_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_001_src3_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src3_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_001_src3_ready                                                                                                 : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_demux_001:src3_ready
	signal width_adapter_002_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_002:out_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                                                   : std_logic;                      -- width_adapter_002:out_valid -> cmd_xbar_mux_003:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_002:out_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal width_adapter_002_src_data                                                                                                    : std_logic_vector(90 downto 0);  -- width_adapter_002:out_data -> cmd_xbar_mux_003:sink0_data
	signal width_adapter_002_src_ready                                                                                                   : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_002:out_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_001_src16_endofpacket                                                                                          : std_logic;                      -- cmd_xbar_demux_001:src16_endofpacket -> width_adapter_003:in_endofpacket
	signal cmd_xbar_demux_001_src16_valid                                                                                                : std_logic;                      -- cmd_xbar_demux_001:src16_valid -> width_adapter_003:in_valid
	signal cmd_xbar_demux_001_src16_startofpacket                                                                                        : std_logic;                      -- cmd_xbar_demux_001:src16_startofpacket -> width_adapter_003:in_startofpacket
	signal cmd_xbar_demux_001_src16_data                                                                                                 : std_logic_vector(108 downto 0); -- cmd_xbar_demux_001:src16_data -> width_adapter_003:in_data
	signal cmd_xbar_demux_001_src16_channel                                                                                              : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_001:src16_channel -> width_adapter_003:in_channel
	signal cmd_xbar_demux_001_src16_ready                                                                                                : std_logic;                      -- width_adapter_003:in_ready -> cmd_xbar_demux_001:src16_ready
	signal width_adapter_003_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_003:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	signal width_adapter_003_src_valid                                                                                                   : std_logic;                      -- width_adapter_003:out_valid -> burst_adapter_002:sink0_valid
	signal width_adapter_003_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_003:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	signal width_adapter_003_src_data                                                                                                    : std_logic_vector(81 downto 0);  -- width_adapter_003:out_data -> burst_adapter_002:sink0_data
	signal width_adapter_003_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_003:out_channel -> burst_adapter_002:sink0_channel
	signal cmd_xbar_demux_002_src0_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> width_adapter_004:in_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> width_adapter_004:in_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> width_adapter_004:in_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                                                  : std_logic_vector(81 downto 0);  -- cmd_xbar_demux_002:src0_data -> width_adapter_004:in_data
	signal cmd_xbar_demux_002_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_002:src0_channel -> width_adapter_004:in_channel
	signal cmd_xbar_demux_002_src0_ready                                                                                                 : std_logic;                      -- width_adapter_004:in_ready -> cmd_xbar_demux_002:src0_ready
	signal width_adapter_004_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_004:out_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal width_adapter_004_src_valid                                                                                                   : std_logic;                      -- width_adapter_004:out_valid -> cmd_xbar_mux_003:sink1_valid
	signal width_adapter_004_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_004:out_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal width_adapter_004_src_data                                                                                                    : std_logic_vector(90 downto 0);  -- width_adapter_004:out_data -> cmd_xbar_mux_003:sink1_data
	signal width_adapter_004_src_ready                                                                                                   : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_004:out_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_003_src0_endofpacket                                                                                           : std_logic;                      -- cmd_xbar_demux_003:src0_endofpacket -> width_adapter_005:in_endofpacket
	signal cmd_xbar_demux_003_src0_valid                                                                                                 : std_logic;                      -- cmd_xbar_demux_003:src0_valid -> width_adapter_005:in_valid
	signal cmd_xbar_demux_003_src0_startofpacket                                                                                         : std_logic;                      -- cmd_xbar_demux_003:src0_startofpacket -> width_adapter_005:in_startofpacket
	signal cmd_xbar_demux_003_src0_data                                                                                                  : std_logic_vector(81 downto 0);  -- cmd_xbar_demux_003:src0_data -> width_adapter_005:in_data
	signal cmd_xbar_demux_003_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- cmd_xbar_demux_003:src0_channel -> width_adapter_005:in_channel
	signal cmd_xbar_demux_003_src0_ready                                                                                                 : std_logic;                      -- width_adapter_005:in_ready -> cmd_xbar_demux_003:src0_ready
	signal width_adapter_005_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_005:out_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	signal width_adapter_005_src_valid                                                                                                   : std_logic;                      -- width_adapter_005:out_valid -> cmd_xbar_mux_003:sink2_valid
	signal width_adapter_005_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_005:out_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	signal width_adapter_005_src_data                                                                                                    : std_logic_vector(90 downto 0);  -- width_adapter_005:out_data -> cmd_xbar_mux_003:sink2_data
	signal width_adapter_005_src_ready                                                                                                   : std_logic;                      -- cmd_xbar_mux_003:sink2_ready -> width_adapter_005:out_ready
	signal width_adapter_005_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_005:out_channel -> cmd_xbar_mux_003:sink2_channel
	signal rsp_xbar_demux_002_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> width_adapter_006:in_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> width_adapter_006:in_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> width_adapter_006:in_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                                                  : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_002:src0_data -> width_adapter_006:in_data
	signal rsp_xbar_demux_002_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_002:src0_channel -> width_adapter_006:in_channel
	signal rsp_xbar_demux_002_src0_ready                                                                                                 : std_logic;                      -- width_adapter_006:in_ready -> rsp_xbar_demux_002:src0_ready
	signal width_adapter_006_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_006:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal width_adapter_006_src_valid                                                                                                   : std_logic;                      -- width_adapter_006:out_valid -> rsp_xbar_mux:sink2_valid
	signal width_adapter_006_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_006:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal width_adapter_006_src_data                                                                                                    : std_logic_vector(108 downto 0); -- width_adapter_006:out_data -> rsp_xbar_mux:sink2_data
	signal width_adapter_006_src_ready                                                                                                   : std_logic;                      -- rsp_xbar_mux:sink2_ready -> width_adapter_006:out_ready
	signal width_adapter_006_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_006:out_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src1_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> width_adapter_007:in_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> width_adapter_007:in_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> width_adapter_007:in_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                                                  : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_002:src1_data -> width_adapter_007:in_data
	signal rsp_xbar_demux_002_src1_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_002:src1_channel -> width_adapter_007:in_channel
	signal rsp_xbar_demux_002_src1_ready                                                                                                 : std_logic;                      -- width_adapter_007:in_ready -> rsp_xbar_demux_002:src1_ready
	signal width_adapter_007_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal width_adapter_007_src_valid                                                                                                   : std_logic;                      -- width_adapter_007:out_valid -> rsp_xbar_mux_001:sink2_valid
	signal width_adapter_007_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal width_adapter_007_src_data                                                                                                    : std_logic_vector(108 downto 0); -- width_adapter_007:out_data -> rsp_xbar_mux_001:sink2_data
	signal width_adapter_007_src_ready                                                                                                   : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> width_adapter_007:out_ready
	signal width_adapter_007_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_007:out_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_003_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> width_adapter_008:in_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> width_adapter_008:in_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> width_adapter_008:in_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                                                  : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_003:src0_data -> width_adapter_008:in_data
	signal rsp_xbar_demux_003_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_003:src0_channel -> width_adapter_008:in_channel
	signal rsp_xbar_demux_003_src0_ready                                                                                                 : std_logic;                      -- width_adapter_008:in_ready -> rsp_xbar_demux_003:src0_ready
	signal width_adapter_008_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal width_adapter_008_src_valid                                                                                                   : std_logic;                      -- width_adapter_008:out_valid -> rsp_xbar_mux_001:sink3_valid
	signal width_adapter_008_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal width_adapter_008_src_data                                                                                                    : std_logic_vector(108 downto 0); -- width_adapter_008:out_data -> rsp_xbar_mux_001:sink3_data
	signal width_adapter_008_src_ready                                                                                                   : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> width_adapter_008:out_ready
	signal width_adapter_008_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_008:out_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> width_adapter_009:in_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> width_adapter_009:in_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> width_adapter_009:in_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                                                  : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_003:src1_data -> width_adapter_009:in_data
	signal rsp_xbar_demux_003_src1_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_003:src1_channel -> width_adapter_009:in_channel
	signal rsp_xbar_demux_003_src1_ready                                                                                                 : std_logic;                      -- width_adapter_009:in_ready -> rsp_xbar_demux_003:src1_ready
	signal width_adapter_009_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_009:out_endofpacket -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal width_adapter_009_src_valid                                                                                                   : std_logic;                      -- width_adapter_009:out_valid -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	signal width_adapter_009_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_009:out_startofpacket -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal width_adapter_009_src_data                                                                                                    : std_logic_vector(81 downto 0);  -- width_adapter_009:out_data -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	signal width_adapter_009_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_009:out_channel -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_003_src2_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_003:src2_endofpacket -> width_adapter_010:in_endofpacket
	signal rsp_xbar_demux_003_src2_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_003:src2_valid -> width_adapter_010:in_valid
	signal rsp_xbar_demux_003_src2_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_003:src2_startofpacket -> width_adapter_010:in_startofpacket
	signal rsp_xbar_demux_003_src2_data                                                                                                  : std_logic_vector(90 downto 0);  -- rsp_xbar_demux_003:src2_data -> width_adapter_010:in_data
	signal rsp_xbar_demux_003_src2_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_003:src2_channel -> width_adapter_010:in_channel
	signal rsp_xbar_demux_003_src2_ready                                                                                                 : std_logic;                      -- width_adapter_010:in_ready -> rsp_xbar_demux_003:src2_ready
	signal width_adapter_010_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_010:out_endofpacket -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal width_adapter_010_src_valid                                                                                                   : std_logic;                      -- width_adapter_010:out_valid -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	signal width_adapter_010_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_010:out_startofpacket -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal width_adapter_010_src_data                                                                                                    : std_logic_vector(81 downto 0);  -- width_adapter_010:out_data -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	signal width_adapter_010_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_010:out_channel -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_016_src0_endofpacket                                                                                           : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> width_adapter_011:in_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                                                 : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> width_adapter_011:in_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                                                         : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> width_adapter_011:in_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                                                  : std_logic_vector(81 downto 0);  -- rsp_xbar_demux_016:src0_data -> width_adapter_011:in_data
	signal rsp_xbar_demux_016_src0_channel                                                                                               : std_logic_vector(16 downto 0);  -- rsp_xbar_demux_016:src0_channel -> width_adapter_011:in_channel
	signal rsp_xbar_demux_016_src0_ready                                                                                                 : std_logic;                      -- width_adapter_011:in_ready -> rsp_xbar_demux_016:src0_ready
	signal width_adapter_011_src_endofpacket                                                                                             : std_logic;                      -- width_adapter_011:out_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	signal width_adapter_011_src_valid                                                                                                   : std_logic;                      -- width_adapter_011:out_valid -> rsp_xbar_mux_001:sink16_valid
	signal width_adapter_011_src_startofpacket                                                                                           : std_logic;                      -- width_adapter_011:out_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	signal width_adapter_011_src_data                                                                                                    : std_logic_vector(108 downto 0); -- width_adapter_011:out_data -> rsp_xbar_mux_001:sink16_data
	signal width_adapter_011_src_ready                                                                                                   : std_logic;                      -- rsp_xbar_mux_001:sink16_ready -> width_adapter_011:out_ready
	signal width_adapter_011_src_channel                                                                                                 : std_logic_vector(16 downto 0);  -- width_adapter_011:out_channel -> rsp_xbar_mux_001:sink16_channel
	signal irq_mapper_receiver0_irq                                                                                                      : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                                                      : std_logic;                      -- timer_system:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                                                      : std_logic;                      -- timer_timestamp:irq -> irq_mapper:receiver2_irq
	signal cpu_d_irq_irq                                                                                                                 : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> CPU:d_irq
	signal reset_n_ports_inv                                                                                                             : std_logic;                      -- reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                                                     : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_write:inv -> sdram_0:az_wr_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv                                                                      : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_read:inv -> sdram_0:az_rd_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                                                : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram_0:az_be_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                                  : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                                   : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal timer_system_s1_translator_avalon_anti_slave_0_write_ports_inv                                                                : std_logic;                      -- timer_system_s1_translator_avalon_anti_slave_0_write:inv -> timer_system:write_n
	signal timer_timestamp_s1_translator_avalon_anti_slave_0_write_ports_inv                                                             : std_logic;                      -- timer_timestamp_s1_translator_avalon_anti_slave_0_write:inv -> timer_timestamp:write_n
	signal red_leds_s1_translator_avalon_anti_slave_0_write_ports_inv                                                                    : std_logic;                      -- red_leds_s1_translator_avalon_anti_slave_0_write:inv -> red_leds:write_n
	signal green_leds_s1_translator_avalon_anti_slave_0_write_ports_inv                                                                  : std_logic;                      -- green_leds_s1_translator_avalon_anti_slave_0_write:inv -> green_leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                                                      : std_logic;                      -- rst_controller_reset_out_reset:inv -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, Barcode_scan_0:avs_s1_reset_n, Barcode_scan_0:reset_n, CPU:reset_n, green_leds:reset_n, jtag_uart_0:rst_n, lcd:reset_n, red_leds:reset_n, sdram_0:reset_n, switch:reset_n, sysid_qsys_0:reset_n, timer_system:reset_n, timer_timestamp:reset_n]
	signal clock_signals_sys_clk_reset_reset_ports_inv                                                                                   : std_logic;                      -- clock_signals_sys_clk_reset_reset:inv -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2]

begin

	onchip_memory : component SOPC_Video_Onchip_Memory
		port map (
			clk        => clock_signals_sys_clk_clk,                                  --   clk1.clk
			address    => onchip_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => onchip_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => onchip_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                          --       .reset_req
		);

	dual_clock_fifo : component SOPC_Video_Dual_Clock_FIFO
		port map (
			clk_stream_in            => clock_signals_sys_clk_clk,                             --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                        --   clock_stream_in_reset.reset
			clk_stream_out           => clock_signals_vga_clk_clk,                             --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,                    --  clock_stream_out_reset.reset
			stream_in_ready          => pixel_rgb_resampler_avalon_rgb_source_ready,           --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => pixel_rgb_resampler_avalon_rgb_source_startofpacket,   --                        .startofpacket
			stream_in_endofpacket    => pixel_rgb_resampler_avalon_rgb_source_endofpacket,     --                        .endofpacket
			stream_in_valid          => pixel_rgb_resampler_avalon_rgb_source_valid,           --                        .valid
			stream_in_data           => pixel_rgb_resampler_avalon_rgb_source_data,            --                        .data
			stream_out_ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	pixel_buffer : component SOPC_Video_Pixel_Buffer
		port map (
			clk           => clock_signals_sys_clk_clk,                                                   --        clock_reset.clk
			reset         => rst_controller_reset_out_reset,                                              --  clock_reset_reset.reset
			SRAM_DQ       => SRAM_DQ_to_and_from_the_Pixel_Buffer,                                        -- external_interface.export
			SRAM_ADDR     => SRAM_ADDR_from_the_Pixel_Buffer,                                             --                   .export
			SRAM_LB_N     => SRAM_LB_N_from_the_Pixel_Buffer,                                             --                   .export
			SRAM_UB_N     => SRAM_UB_N_from_the_Pixel_Buffer,                                             --                   .export
			SRAM_CE_N     => SRAM_CE_N_from_the_Pixel_Buffer,                                             --                   .export
			SRAM_OE_N     => SRAM_OE_N_from_the_Pixel_Buffer,                                             --                   .export
			SRAM_WE_N     => SRAM_WE_N_from_the_Pixel_Buffer,                                             --                   .export
			address       => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address,       --  avalon_sram_slave.address
			byteenable    => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,    --                   .byteenable
			read          => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read,          --                   .read
			write         => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write,         --                   .write
			writedata     => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,     --                   .writedata
			readdata      => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,      --                   .readdata
			readdatavalid => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid  --                   .readdatavalid
		);

	pixel_buffer_dma : component SOPC_Video_Pixel_Buffer_DMA
		port map (
			clk                  => clock_signals_sys_clk_clk,                                                       --             clock_reset.clk
			reset                => rst_controller_reset_out_reset,                                                  --       clock_reset_reset.reset
			master_readdatavalid => pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,                          -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,                            --                        .waitrequest
			master_address       => pixel_buffer_dma_avalon_pixel_dma_master_address,                                --                        .address
			master_arbiterlock   => pixel_buffer_dma_avalon_pixel_dma_master_lock,                                   --                        .lock
			master_read          => pixel_buffer_dma_avalon_pixel_dma_master_read,                                   --                        .read
			master_readdata      => pixel_buffer_dma_avalon_pixel_dma_master_readdata,                               --                        .readdata
			slave_address        => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address,    --    avalon_control_slave.address
			slave_byteenable     => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable, --                        .byteenable
			slave_read           => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read,       --                        .read
			slave_write          => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write,      --                        .write
			slave_writedata      => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata,  --                        .writedata
			slave_readdata       => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata,   --                        .readdata
			stream_ready         => pixel_buffer_dma_avalon_pixel_source_ready,                                      --     avalon_pixel_source.ready
			stream_startofpacket => pixel_buffer_dma_avalon_pixel_source_startofpacket,                              --                        .startofpacket
			stream_endofpacket   => pixel_buffer_dma_avalon_pixel_source_endofpacket,                                --                        .endofpacket
			stream_valid         => pixel_buffer_dma_avalon_pixel_source_valid,                                      --                        .valid
			stream_data          => pixel_buffer_dma_avalon_pixel_source_data                                        --                        .data
		);

	pixel_rgb_resampler : component SOPC_Video_Pixel_RGB_Resampler
		port map (
			clk                      => clock_signals_sys_clk_clk,                           --       clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                      -- clock_reset_reset.reset
			stream_in_startofpacket  => pixel_buffer_dma_avalon_pixel_source_startofpacket,  --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => pixel_buffer_dma_avalon_pixel_source_endofpacket,    --                  .endofpacket
			stream_in_valid          => pixel_buffer_dma_avalon_pixel_source_valid,          --                  .valid
			stream_in_ready          => pixel_buffer_dma_avalon_pixel_source_ready,          --                  .ready
			stream_in_data           => pixel_buffer_dma_avalon_pixel_source_data,           --                  .data
			stream_out_ready         => pixel_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => pixel_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => pixel_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => pixel_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => pixel_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	vga_controller : component SOPC_Video_VGA_Controller
		port map (
			clk           => clock_signals_vga_clk_clk,                             --        clock_reset.clk
			reset         => rst_controller_001_reset_out_reset,                    --  clock_reset_reset.reset
			data          => dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => VGA_CLK_from_the_VGA_Controller,                       -- external_interface.export
			VGA_HS        => VGA_HS_from_the_VGA_Controller,                        --                   .export
			VGA_VS        => VGA_VS_from_the_VGA_Controller,                        --                   .export
			VGA_BLANK     => VGA_BLANK_from_the_VGA_Controller,                     --                   .export
			VGA_SYNC      => VGA_SYNC_from_the_VGA_Controller,                      --                   .export
			VGA_R         => VGA_R_from_the_VGA_Controller,                         --                   .export
			VGA_G         => VGA_G_from_the_VGA_Controller,                         --                   .export
			VGA_B         => VGA_B_from_the_VGA_Controller                          --                   .export
		);

	video_in_decoder : component SOPC_Video_Video_In_Decoder
		port map (
			clk                      => clock_signals_sys_clk_clk,                            --           clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                       --     clock_reset_reset.reset
			stream_out_ready         => video_in_decoder_avalon_decoder_source_ready,         -- avalon_decoder_source.ready
			stream_out_startofpacket => video_in_decoder_avalon_decoder_source_startofpacket, --                      .startofpacket
			stream_out_endofpacket   => video_in_decoder_avalon_decoder_source_endofpacket,   --                      .endofpacket
			stream_out_valid         => video_in_decoder_avalon_decoder_source_valid,         --                      .valid
			stream_out_data          => video_in_decoder_avalon_decoder_source_data,          --                      .data
			PIXEL_CLK                => Video_In_Decoder_external_interface_PIXEL_CLK,        --    external_interface.export
			LINE_VALID               => Video_In_Decoder_external_interface_LINE_VALID,       --                      .export
			FRAME_VALID              => Video_In_Decoder_external_interface_FRAME_VALID,      --                      .export
			pixel_clk_reset          => Video_In_Decoder_external_interface_pixel_clk_reset,  --                      .export
			PIXEL_DATA               => Video_In_Decoder_external_interface_PIXEL_DATA        --                      .export
		);

	video_dma : component SOPC_Video_Video_DMA
		port map (
			clk                  => clock_signals_sys_clk_clk,                                                    --              clock_reset.clk
			reset                => rst_controller_reset_out_reset,                                               --        clock_reset_reset.reset
			stream_data          => barcode_scan_0_avalon_streaming_source_data,                                  --          avalon_dma_sink.data
			stream_startofpacket => barcode_scan_0_avalon_streaming_source_startofpacket,                         --                         .startofpacket
			stream_endofpacket   => barcode_scan_0_avalon_streaming_source_endofpacket,                           --                         .endofpacket
			stream_valid         => barcode_scan_0_avalon_streaming_source_valid,                                 --                         .valid
			stream_ready         => barcode_scan_0_avalon_streaming_source_ready,                                 --                         .ready
			slave_address        => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable, --                         .byteenable
			slave_read           => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read,       --                         .read
			slave_write          => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write,      --                         .write
			slave_writedata      => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata,  --                         .writedata
			slave_readdata       => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata,   --                         .readdata
			master_address       => video_dma_avalon_dma_master_address,                                          --        avalon_dma_master.address
			master_waitrequest   => video_dma_avalon_dma_master_waitrequest,                                      --                         .waitrequest
			master_write         => video_dma_avalon_dma_master_write,                                            --                         .write
			master_writedata     => video_dma_avalon_dma_master_writedata                                         --                         .writedata
		);

	av_config : component SOPC_Video_AV_Config
		port map (
			clk         => clock_signals_sys_clk_clk,                                                   --            clock_reset.clk
			reset       => rst_controller_reset_out_reset,                                              --      clock_reset_reset.reset
			address     => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address,     -- avalon_av_config_slave.address
			byteenable  => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable,  --                       .byteenable
			read        => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read,        --                       .read
			write       => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write,       --                       .write
			writedata   => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata,   --                       .writedata
			readdata    => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata,    --                       .readdata
			waitrequest => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest, --                       .waitrequest
			I2C_SDAT    => I2C_SDAT_to_and_from_the_AV_Config,                                          --     external_interface.export
			I2C_SCLK    => I2C_SCLK_from_the_AV_Config                                                  --                       .export
		);

	cpu : component SOPC_Video_CPU
		port map (
			clk                                   => clock_signals_sys_clk_clk,                                        --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			E_ci_multi_done                       => cpu_custom_instruction_master_done,                               -- custom_instruction_master.done
			E_ci_multi_clk_en                     => cpu_custom_instruction_master_clk_en,                             --                          .clk_en
			E_ci_multi_start                      => cpu_custom_instruction_master_start,                              --                          .start
			E_ci_result                           => cpu_custom_instruction_master_result,                             --                          .result
			D_ci_a                                => cpu_custom_instruction_master_a,                                  --                          .a
			D_ci_b                                => cpu_custom_instruction_master_b,                                  --                          .b
			D_ci_c                                => cpu_custom_instruction_master_c,                                  --                          .c
			D_ci_n                                => cpu_custom_instruction_master_n,                                  --                          .n
			D_ci_readra                           => cpu_custom_instruction_master_readra,                             --                          .readra
			D_ci_readrb                           => cpu_custom_instruction_master_readrb,                             --                          .readrb
			D_ci_writerc                          => cpu_custom_instruction_master_writerc,                            --                          .writerc
			E_ci_dataa                            => cpu_custom_instruction_master_dataa,                              --                          .dataa
			E_ci_datab                            => cpu_custom_instruction_master_datab,                              --                          .datab
			E_ci_multi_clock                      => cpu_custom_instruction_master_clk,                                --                          .clk
			E_ci_multi_reset                      => cpu_custom_instruction_master_reset,                              --                          .reset
			W_ci_estatus                          => cpu_custom_instruction_master_estatus,                            --                          .estatus
			W_ci_ipending                         => cpu_custom_instruction_master_ipending                            --                          .ipending
		);

	clock_signals : component SOPC_Video_Clock_Signals
		port map (
			CLOCK_50    => clk_0,                              --       clk_in_primary.clk
			reset       => rst_controller_002_reset_out_reset, -- clk_in_primary_reset.reset
			sys_clk     => clock_signals_sys_clk_clk,          --              sys_clk.clk
			sys_reset_n => clock_signals_sys_clk_reset_reset,  --        sys_clk_reset.reset_n
			SDRAM_CLK   => sdram_clk_clk,                      --            sdram_clk.clk
			VGA_CLK     => clock_signals_vga_clk_clk           --              vga_clk.clk
		);

	jtag_uart_0 : component SOPC_Video_jtag_uart_0
		port map (
			clk            => clock_signals_sys_clk_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                     --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                      --               irq.irq
		);

	video_bayer_resampler : component SOPC_Video_video_bayer_resampler
		port map (
			clk                      => clock_signals_sys_clk_clk,                               --         clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                          --   clock_reset_reset.reset
			stream_in_data           => video_in_decoder_avalon_decoder_source_data,             --   avalon_bayer_sink.data
			stream_in_startofpacket  => video_in_decoder_avalon_decoder_source_startofpacket,    --                    .startofpacket
			stream_in_endofpacket    => video_in_decoder_avalon_decoder_source_endofpacket,      --                    .endofpacket
			stream_in_valid          => video_in_decoder_avalon_decoder_source_valid,            --                    .valid
			stream_in_ready          => video_in_decoder_avalon_decoder_source_ready,            --                    .ready
			stream_out_ready         => video_bayer_resampler_avalon_bayer_source_ready,         -- avalon_bayer_source.ready
			stream_out_data          => video_bayer_resampler_avalon_bayer_source_data,          --                    .data
			stream_out_startofpacket => video_bayer_resampler_avalon_bayer_source_startofpacket, --                    .startofpacket
			stream_out_endofpacket   => video_bayer_resampler_avalon_bayer_source_endofpacket,   --                    .endofpacket
			stream_out_valid         => video_bayer_resampler_avalon_bayer_source_valid          --                    .valid
		);

	video_clipper_0 : component SOPC_Video_video_clipper_0
		port map (
			clk                      => clock_signals_sys_clk_clk,                               --           clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                          --     clock_reset_reset.reset
			stream_in_data           => video_bayer_resampler_avalon_bayer_source_data,          --   avalon_clipper_sink.data
			stream_in_startofpacket  => video_bayer_resampler_avalon_bayer_source_startofpacket, --                      .startofpacket
			stream_in_endofpacket    => video_bayer_resampler_avalon_bayer_source_endofpacket,   --                      .endofpacket
			stream_in_valid          => video_bayer_resampler_avalon_bayer_source_valid,         --                      .valid
			stream_in_ready          => video_bayer_resampler_avalon_bayer_source_ready,         --                      .ready
			stream_out_ready         => video_clipper_0_avalon_clipper_source_ready,             -- avalon_clipper_source.ready
			stream_out_data          => video_clipper_0_avalon_clipper_source_data,              --                      .data
			stream_out_startofpacket => video_clipper_0_avalon_clipper_source_startofpacket,     --                      .startofpacket
			stream_out_endofpacket   => video_clipper_0_avalon_clipper_source_endofpacket,       --                      .endofpacket
			stream_out_valid         => video_clipper_0_avalon_clipper_source_valid              --                      .valid
		);

	video_scaler_0 : component SOPC_Video_video_scaler_0
		port map (
			clk                      => clock_signals_sys_clk_clk,                           --          clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                      --    clock_reset_reset.reset
			stream_in_startofpacket  => video_clipper_0_avalon_clipper_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_clipper_0_avalon_clipper_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_clipper_0_avalon_clipper_source_valid,         --                     .valid
			stream_in_ready          => video_clipper_0_avalon_clipper_source_ready,         --                     .ready
			stream_in_data           => video_clipper_0_avalon_clipper_source_data,          --                     .data
			stream_out_ready         => video_scaler_0_avalon_scaler_source_ready,           -- avalon_scaler_source.ready
			stream_out_startofpacket => video_scaler_0_avalon_scaler_source_startofpacket,   --                     .startofpacket
			stream_out_endofpacket   => video_scaler_0_avalon_scaler_source_endofpacket,     --                     .endofpacket
			stream_out_valid         => video_scaler_0_avalon_scaler_source_valid,           --                     .valid
			stream_out_data          => video_scaler_0_avalon_scaler_source_data             --                     .data
		);

	video_rgb_resampler_0 : component SOPC_Video_video_rgb_resampler_0
		port map (
			clk                      => clock_signals_sys_clk_clk,                             --       clock_reset.clk
			reset                    => rst_controller_reset_out_reset,                        -- clock_reset_reset.reset
			stream_in_startofpacket  => video_scaler_0_avalon_scaler_source_startofpacket,     --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_scaler_0_avalon_scaler_source_endofpacket,       --                  .endofpacket
			stream_in_valid          => video_scaler_0_avalon_scaler_source_valid,             --                  .valid
			stream_in_ready          => video_scaler_0_avalon_scaler_source_ready,             --                  .ready
			stream_in_data           => video_scaler_0_avalon_scaler_source_data,              --                  .data
			stream_out_ready         => video_rgb_resampler_0_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => video_rgb_resampler_0_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_rgb_resampler_0_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_rgb_resampler_0_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => video_rgb_resampler_0_avalon_rgb_source_data           --                  .data
		);

	sysid_qsys_0 : component SOPC_Video_sysid_qsys_0
		port map (
			clock    => clock_signals_sys_clk_clk,                                            --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                             --         reset.reset_n
			readdata => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	sdram_0 : component SOPC_Video_sdram_0
		port map (
			clk            => clock_signals_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                       -- reset.reset_n
			az_addr        => sdram_0_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_0_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_0_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                                --  wire.export
			zs_ba          => sdram_wire_ba,                                                  --      .export
			zs_cas_n       => sdram_wire_cas_n,                                               --      .export
			zs_cke         => sdram_wire_cke,                                                 --      .export
			zs_cs_n        => sdram_wire_cs_n,                                                --      .export
			zs_dq          => sdram_wire_dq,                                                  --      .export
			zs_dqm         => sdram_wire_dqm,                                                 --      .export
			zs_ras_n       => sdram_wire_ras_n,                                               --      .export
			zs_we_n        => sdram_wire_we_n                                                 --      .export
		);

	timer_system : component SOPC_Video_timer_system
		port map (
			clk        => clock_signals_sys_clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                       -- reset.reset_n
			address    => timer_system_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_system_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_system_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_system_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_system_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                        --   irq.irq
		);

	timer_timestamp : component SOPC_Video_timer_system
		port map (
			clk        => clock_signals_sys_clk_clk,                                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                          -- reset.reset_n
			address    => timer_timestamp_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_timestamp_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_timestamp_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_timestamp_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                                           --   irq.irq
		);

	lcd : component SOPC_Video_lcd
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,                       --         reset.reset_n
			clk           => clock_signals_sys_clk_clk,                                      --           clk.clk
			begintransfer => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer, -- control_slave.begintransfer
			read          => lcd_control_slave_translator_avalon_anti_slave_0_read,          --              .read
			write         => lcd_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			readdata      => lcd_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			writedata     => lcd_control_slave_translator_avalon_anti_slave_0_writedata,     --              .writedata
			address       => lcd_control_slave_translator_avalon_anti_slave_0_address,       --              .address
			LCD_RS        => lcd_ext_RS,                                                     --      external.export
			LCD_RW        => lcd_ext_RW,                                                     --              .export
			LCD_data      => lcd_ext_data,                                                   --              .export
			LCD_E         => lcd_ext_E                                                       --              .export
		);

	red_leds : component SOPC_Video_red_leds
		port map (
			clk        => clock_signals_sys_clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => red_leds_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => red_leds_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => red_leds_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => red_leds_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => red_leds_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => red_leds_ext_export                                         -- external_connection.export
		);

	green_leds : component SOPC_Video_red_leds
		port map (
			clk        => clock_signals_sys_clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => green_leds_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => green_leds_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => green_leds_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => green_leds_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => green_leds_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => green_leds_ext_export                                         -- external_connection.export
		);

	switch : component SOPC_Video_switch
		port map (
			clk      => clock_signals_sys_clk_clk,                         --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => switch_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => switch_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => switch_ext_export                                  -- external_connection.export
		);

	nios_custom_instr_floating_point_0 : component fpoint_wrapper
		generic map (
			useDivider => 0
		)
		port map (
			clk    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- s1.clk
			clk_en => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --   .clk_en
			dataa  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --   .dataa
			datab  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --   .datab
			n      => cpu_custom_instruction_master_multi_slave_translator0_ci_master_n,      --   .n
			reset  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --   .reset
			start  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --   .start
			done   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done,   --   .done
			result => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result  --   .result
		);

	altera_up_sd_card_avalon_interface_0 : component Altera_UP_SD_Card_Avalon_Interface
		port map (
			i_avalon_chip_select => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect,  -- avalon_sdcard_slave.chipselect
			i_avalon_address     => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address,     --                    .address
			i_avalon_read        => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read,        --                    .read
			i_avalon_write       => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write,       --                    .write
			i_avalon_byteenable  => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable,  --                    .byteenable
			i_avalon_writedata   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata,   --                    .writedata
			o_avalon_readdata    => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata,    --                    .readdata
			o_avalon_waitrequest => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest, --                    .waitrequest
			i_clock              => clock_signals_sys_clk_clk,                                                                           --          clock_sink.clk
			i_reset_n            => rst_controller_reset_out_reset_ports_inv,                                                            --    clock_sink_reset.reset_n
			b_SD_cmd             => altera_up_sd_card_b_SD_cmd,                                                                          --         conduit_end.export
			b_SD_dat             => altera_up_sd_card_b_SD_dat,                                                                          --                    .export
			b_SD_dat3            => altera_up_sd_card_b_SD_dat3,                                                                         --                    .export
			o_SD_clock           => altera_up_sd_card_o_SD_clock                                                                         --                    .export
		);

	barcode_scan_0 : component pixel_scan
		port map (
			avs_s1_write             => barcode_scan_0_s1_translator_avalon_anti_slave_0_write,      --                      s1.write
			avs_s1_read              => barcode_scan_0_s1_translator_avalon_anti_slave_0_read,       --                        .read
			avs_s1_chipselect        => barcode_scan_0_s1_translator_avalon_anti_slave_0_chipselect, --                        .chipselect
			avs_s1_address           => barcode_scan_0_s1_translator_avalon_anti_slave_0_address,    --                        .address
			avs_s1_writedata         => barcode_scan_0_s1_translator_avalon_anti_slave_0_writedata,  --                        .writedata
			avs_s1_readdata          => barcode_scan_0_s1_translator_avalon_anti_slave_0_readdata,   --                        .readdata
			ast_sink_ready           => video_rgb_resampler_0_avalon_rgb_source_ready,               --   avalon_streaming_sink.ready
			ast_sink_valid           => video_rgb_resampler_0_avalon_rgb_source_valid,               --                        .valid
			ast_sink_startofpacket   => video_rgb_resampler_0_avalon_rgb_source_startofpacket,       --                        .startofpacket
			ast_sink_endofpacket     => video_rgb_resampler_0_avalon_rgb_source_endofpacket,         --                        .endofpacket
			ast_sink_data            => video_rgb_resampler_0_avalon_rgb_source_data,                --                        .data
			clk                      => clock_signals_sys_clk_clk,                                   --                clock_st.clk
			reset_n                  => rst_controller_reset_out_reset_ports_inv,                    --                reset_st.reset_n
			avs_s1_clk               => clock_signals_sys_clk_clk,                                   --                clock_mm.clk
			avs_s1_reset_n           => rst_controller_reset_out_reset_ports_inv,                    --                reset_mm.reset_n
			ast_source_valid         => barcode_scan_0_avalon_streaming_source_valid,                -- avalon_streaming_source.valid
			ast_source_endofpacket   => barcode_scan_0_avalon_streaming_source_endofpacket,          --                        .endofpacket
			ast_source_data          => barcode_scan_0_avalon_streaming_source_data,                 --                        .data
			ast_source_startofpacket => barcode_scan_0_avalon_streaming_source_startofpacket,        --                        .startofpacket
			ast_source_ready         => barcode_scan_0_avalon_streaming_source_ready,                --                        .ready
			debug_state              => debug_export,                                                --                   debug.export
			restart                  => restart_export                                               --                 restart.export
		);

	cpu_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa          => cpu_custom_instruction_master_dataa,                              --        ci_slave.dataa
			ci_slave_datab          => cpu_custom_instruction_master_datab,                              --                .datab
			ci_slave_result         => cpu_custom_instruction_master_result,                             --                .result
			ci_slave_n              => cpu_custom_instruction_master_n,                                  --                .n
			ci_slave_readra         => cpu_custom_instruction_master_readra,                             --                .readra
			ci_slave_readrb         => cpu_custom_instruction_master_readrb,                             --                .readrb
			ci_slave_writerc        => cpu_custom_instruction_master_writerc,                            --                .writerc
			ci_slave_a              => cpu_custom_instruction_master_a,                                  --                .a
			ci_slave_b              => cpu_custom_instruction_master_b,                                  --                .b
			ci_slave_c              => cpu_custom_instruction_master_c,                                  --                .c
			ci_slave_ipending       => cpu_custom_instruction_master_ipending,                           --                .ipending
			ci_slave_estatus        => cpu_custom_instruction_master_estatus,                            --                .estatus
			ci_slave_multi_clk      => cpu_custom_instruction_master_clk,                                --                .clk
			ci_slave_multi_reset    => cpu_custom_instruction_master_reset,                              --                .reset
			ci_slave_multi_clken    => cpu_custom_instruction_master_clk_en,                             --                .clk_en
			ci_slave_multi_start    => cpu_custom_instruction_master_start,                              --                .start
			ci_slave_multi_done     => cpu_custom_instruction_master_done,                               --                .done
			comb_ci_master_dataa    => open,                                                             --  comb_ci_master.dataa
			comb_ci_master_datab    => open,                                                             --                .datab
			comb_ci_master_result   => open,                                                             --                .result
			comb_ci_master_n        => open,                                                             --                .n
			comb_ci_master_readra   => open,                                                             --                .readra
			comb_ci_master_readrb   => open,                                                             --                .readrb
			comb_ci_master_writerc  => open,                                                             --                .writerc
			comb_ci_master_a        => open,                                                             --                .a
			comb_ci_master_b        => open,                                                             --                .b
			comb_ci_master_c        => open,                                                             --                .c
			comb_ci_master_ipending => open,                                                             --                .ipending
			comb_ci_master_estatus  => open,                                                             --                .estatus
			multi_ci_master_clk     => cpu_custom_instruction_master_translator_multi_ci_master_clk,     -- multi_ci_master.clk
			multi_ci_master_reset   => cpu_custom_instruction_master_translator_multi_ci_master_reset,   --                .reset
			multi_ci_master_clken   => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,  --                .clk_en
			multi_ci_master_start   => cpu_custom_instruction_master_translator_multi_ci_master_start,   --                .start
			multi_ci_master_done    => cpu_custom_instruction_master_translator_multi_ci_master_done,    --                .done
			multi_ci_master_dataa   => cpu_custom_instruction_master_translator_multi_ci_master_dataa,   --                .dataa
			multi_ci_master_datab   => cpu_custom_instruction_master_translator_multi_ci_master_datab,   --                .datab
			multi_ci_master_result  => cpu_custom_instruction_master_translator_multi_ci_master_result,  --                .result
			multi_ci_master_n       => cpu_custom_instruction_master_translator_multi_ci_master_n,       --                .n
			multi_ci_master_readra  => cpu_custom_instruction_master_translator_multi_ci_master_readra,  --                .readra
			multi_ci_master_readrb  => cpu_custom_instruction_master_translator_multi_ci_master_readrb,  --                .readrb
			multi_ci_master_writerc => cpu_custom_instruction_master_translator_multi_ci_master_writerc, --                .writerc
			multi_ci_master_a       => cpu_custom_instruction_master_translator_multi_ci_master_a,       --                .a
			multi_ci_master_b       => cpu_custom_instruction_master_translator_multi_ci_master_b,       --                .b
			multi_ci_master_c       => cpu_custom_instruction_master_translator_multi_ci_master_c,       --                .c
			ci_slave_multi_dataa    => "00000000000000000000000000000000",                               --     (terminated)
			ci_slave_multi_datab    => "00000000000000000000000000000000",                               --     (terminated)
			ci_slave_multi_result   => open,                                                             --     (terminated)
			ci_slave_multi_n        => "00000000",                                                       --     (terminated)
			ci_slave_multi_readra   => '0',                                                              --     (terminated)
			ci_slave_multi_readrb   => '0',                                                              --     (terminated)
			ci_slave_multi_writerc  => '0',                                                              --     (terminated)
			ci_slave_multi_a        => "00000",                                                          --     (terminated)
			ci_slave_multi_b        => "00000",                                                          --     (terminated)
			ci_slave_multi_c        => "00000"                                                           --     (terminated)
		);

	cpu_custom_instruction_master_multi_xconnect : component SOPC_Video_CPU_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa      => cpu_custom_instruction_master_translator_multi_ci_master_dataa,   --   ci_slave.dataa
			ci_slave_datab      => cpu_custom_instruction_master_translator_multi_ci_master_datab,   --           .datab
			ci_slave_result     => cpu_custom_instruction_master_translator_multi_ci_master_result,  --           .result
			ci_slave_n          => cpu_custom_instruction_master_translator_multi_ci_master_n,       --           .n
			ci_slave_readra     => cpu_custom_instruction_master_translator_multi_ci_master_readra,  --           .readra
			ci_slave_readrb     => cpu_custom_instruction_master_translator_multi_ci_master_readrb,  --           .readrb
			ci_slave_writerc    => cpu_custom_instruction_master_translator_multi_ci_master_writerc, --           .writerc
			ci_slave_a          => cpu_custom_instruction_master_translator_multi_ci_master_a,       --           .a
			ci_slave_b          => cpu_custom_instruction_master_translator_multi_ci_master_b,       --           .b
			ci_slave_c          => cpu_custom_instruction_master_translator_multi_ci_master_c,       --           .c
			ci_slave_ipending   => open,                                                             --           .ipending
			ci_slave_estatus    => open,                                                             --           .estatus
			ci_slave_clk        => cpu_custom_instruction_master_translator_multi_ci_master_clk,     --           .clk
			ci_slave_reset      => cpu_custom_instruction_master_translator_multi_ci_master_reset,   --           .reset
			ci_slave_clken      => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,  --           .clk_en
			ci_slave_start      => cpu_custom_instruction_master_translator_multi_ci_master_start,   --           .start
			ci_slave_done       => cpu_custom_instruction_master_translator_multi_ci_master_done,    --           .done
			ci_master0_dataa    => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,    -- ci_master0.dataa
			ci_master0_datab    => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,    --           .datab
			ci_master0_result   => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,   --           .result
			ci_master0_n        => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,        --           .n
			ci_master0_readra   => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,   --           .readra
			ci_master0_readrb   => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,   --           .readrb
			ci_master0_writerc  => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,  --           .writerc
			ci_master0_a        => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,        --           .a
			ci_master0_b        => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,        --           .b
			ci_master0_c        => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,        --           .c
			ci_master0_ipending => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending, --           .ipending
			ci_master0_estatus  => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,  --           .estatus
			ci_master0_clk      => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,      --           .clk
			ci_master0_reset    => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,    --           .reset
			ci_master0_clken    => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,   --           .clk_en
			ci_master0_start    => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,    --           .start
			ci_master0_done     => cpu_custom_instruction_master_multi_xconnect_ci_master0_done      --           .done
		);

	cpu_custom_instruction_master_multi_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 2,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa     => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab     => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result    => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n         => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc   => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a         => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b         => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c         => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending  => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus   => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk       => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken     => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset     => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start     => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done      => cpu_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_n        => cpu_custom_instruction_master_multi_slave_translator0_ci_master_n,      --          .n
			ci_master_clk      => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_readra   => open,                                                                   -- (terminated)
			ci_master_readrb   => open,                                                                   -- (terminated)
			ci_master_writerc  => open,                                                                   -- (terminated)
			ci_master_a        => open,                                                                   -- (terminated)
			ci_master_b        => open,                                                                   -- (terminated)
			ci_master_c        => open,                                                                   -- (terminated)
			ci_master_ipending => open,                                                                   -- (terminated)
			ci_master_estatus  => open                                                                    -- (terminated)
		);

	cpu_instruction_master_translator : component sopc_video_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                 --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_readdatavalid         => open,                                                                      --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	cpu_data_master_translator : component sopc_video_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                          --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	pixel_buffer_dma_avalon_pixel_dma_master_translator : component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 8,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 1,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 1,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 1,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                     reset.reset
			uav_address              => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => pixel_buffer_dma_avalon_pixel_dma_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,                                        --                          .waitrequest
			av_read                  => pixel_buffer_dma_avalon_pixel_dma_master_read,                                               --                          .read
			av_readdata              => pixel_buffer_dma_avalon_pixel_dma_master_readdata,                                           --                          .readdata
			av_readdatavalid         => pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,                                      --                          .readdatavalid
			av_lock                  => pixel_buffer_dma_avalon_pixel_dma_master_lock,                                               --                          .lock
			av_burstcount            => "1",                                                                                         --               (terminated)
			av_byteenable            => "1",                                                                                         --               (terminated)
			av_beginbursttransfer    => '0',                                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                                         --               (terminated)
			av_chipselect            => '0',                                                                                         --               (terminated)
			av_write                 => '0',                                                                                         --               (terminated)
			av_writedata             => "00000000",                                                                                  --               (terminated)
			av_debugaccess           => '0',                                                                                         --               (terminated)
			uav_clken                => open,                                                                                        --               (terminated)
			av_clken                 => '1',                                                                                         --               (terminated)
			uav_response             => "00",                                                                                        --               (terminated)
			av_response              => open,                                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                                         --               (terminated)
		);

	video_dma_avalon_dma_master_translator : component sopc_video_video_dma_avalon_dma_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 8,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 1,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 1,
			USE_READ                    => 0,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 1,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                      --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                     reset.reset
			uav_address              => video_dma_avalon_dma_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => video_dma_avalon_dma_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => video_dma_avalon_dma_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => video_dma_avalon_dma_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => video_dma_avalon_dma_master_waitrequest,                                        --                          .waitrequest
			av_write                 => video_dma_avalon_dma_master_write,                                              --                          .write
			av_writedata             => video_dma_avalon_dma_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                            --               (terminated)
			av_byteenable            => "1",                                                                            --               (terminated)
			av_beginbursttransfer    => '0',                                                                            --               (terminated)
			av_begintransfer         => '0',                                                                            --               (terminated)
			av_chipselect            => '0',                                                                            --               (terminated)
			av_read                  => '0',                                                                            --               (terminated)
			av_readdata              => open,                                                                           --               (terminated)
			av_readdatavalid         => open,                                                                           --               (terminated)
			av_lock                  => '0',                                                                            --               (terminated)
			av_debugaccess           => '0',                                                                            --               (terminated)
			uav_clken                => open,                                                                           --               (terminated)
			av_clken                 => '1',                                                                            --               (terminated)
			uav_response             => "00",                                                                           --               (terminated)
			av_response              => open,                                                                           --               (terminated)
			uav_writeresponserequest => open,                                                                           --               (terminated)
			uav_writeresponsevalid   => '0',                                                                            --               (terminated)
			av_writeresponserequest  => '0',                                                                            --               (terminated)
			av_writeresponsevalid    => open                                                                            --               (terminated)
		);

	cpu_jtag_debug_module_translator : component sopc_video_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	onchip_memory_s1_translator : component sopc_video_onchip_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 12,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => onchip_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => onchip_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => onchip_memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	sdram_0_s1_translator : component sopc_video_sdram_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pixel_buffer_avalon_sram_slave_translator : component sopc_video_pixel_buffer_avalon_sram_slave_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                 --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	av_config_avalon_av_config_slave_translator : component sopc_video_av_config_avalon_av_config_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                    reset.reset
			uav_address              => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                                        --              (terminated)
			av_burstcount            => open,                                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                                        --              (terminated)
			av_lock                  => open,                                                                                        --              (terminated)
			av_chipselect            => open,                                                                                        --              (terminated)
			av_clken                 => open,                                                                                        --              (terminated)
			uav_clken                => '0',                                                                                         --              (terminated)
			av_debugaccess           => open,                                                                                        --              (terminated)
			av_outputenable          => open,                                                                                        --              (terminated)
			uav_response             => open,                                                                                        --              (terminated)
			av_response              => "00",                                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                                          --              (terminated)
		);

	video_dma_avalon_dma_control_slave_translator : component sopc_video_video_dma_avalon_dma_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                                --                    reset.reset
			uav_address              => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_begintransfer         => open,                                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                                          --              (terminated)
			av_burstcount            => open,                                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                                          --              (terminated)
			av_lock                  => open,                                                                                          --              (terminated)
			av_chipselect            => open,                                                                                          --              (terminated)
			av_clken                 => open,                                                                                          --              (terminated)
			uav_clken                => '0',                                                                                           --              (terminated)
			av_debugaccess           => open,                                                                                          --              (terminated)
			av_outputenable          => open,                                                                                          --              (terminated)
			uav_response             => open,                                                                                          --              (terminated)
			av_response              => "00",                                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                                            --              (terminated)
		);

	pixel_buffer_dma_avalon_control_slave_translator : component sopc_video_video_dma_avalon_dma_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                                   --                    reset.reset
			uav_address              => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_begintransfer         => open,                                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                                             --              (terminated)
			av_burstcount            => open,                                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                                             --              (terminated)
			av_lock                  => open,                                                                                             --              (terminated)
			av_chipselect            => open,                                                                                             --              (terminated)
			av_clken                 => open,                                                                                             --              (terminated)
			uav_clken                => '0',                                                                                              --              (terminated)
			av_debugaccess           => open,                                                                                             --              (terminated)
			av_outputenable          => open,                                                                                             --              (terminated)
			uav_response             => open,                                                                                             --              (terminated)
			av_response              => "00",                                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                                               --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component sopc_video_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	sysid_qsys_0_control_slave_translator : component sopc_video_sysid_qsys_0_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                        --                    reset.reset
			uav_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                                  --              (terminated)
			av_read                  => open,                                                                                  --              (terminated)
			av_writedata             => open,                                                                                  --              (terminated)
			av_begintransfer         => open,                                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                                  --              (terminated)
			av_burstcount            => open,                                                                                  --              (terminated)
			av_byteenable            => open,                                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                                  --              (terminated)
			av_lock                  => open,                                                                                  --              (terminated)
			av_chipselect            => open,                                                                                  --              (terminated)
			av_clken                 => open,                                                                                  --              (terminated)
			uav_clken                => '0',                                                                                   --              (terminated)
			av_debugaccess           => open,                                                                                  --              (terminated)
			av_outputenable          => open,                                                                                  --              (terminated)
			uav_response             => open,                                                                                  --              (terminated)
			av_response              => "00",                                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                                    --              (terminated)
		);

	timer_system_s1_translator : component sopc_video_timer_system_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                             --                    reset.reset
			uav_address              => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_system_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_system_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_system_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_system_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_system_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                       --              (terminated)
			av_begintransfer         => open,                                                                       --              (terminated)
			av_beginbursttransfer    => open,                                                                       --              (terminated)
			av_burstcount            => open,                                                                       --              (terminated)
			av_byteenable            => open,                                                                       --              (terminated)
			av_readdatavalid         => '0',                                                                        --              (terminated)
			av_waitrequest           => '0',                                                                        --              (terminated)
			av_writebyteenable       => open,                                                                       --              (terminated)
			av_lock                  => open,                                                                       --              (terminated)
			av_clken                 => open,                                                                       --              (terminated)
			uav_clken                => '0',                                                                        --              (terminated)
			av_debugaccess           => open,                                                                       --              (terminated)
			av_outputenable          => open,                                                                       --              (terminated)
			uav_response             => open,                                                                       --              (terminated)
			av_response              => "00",                                                                       --              (terminated)
			uav_writeresponserequest => '0',                                                                        --              (terminated)
			uav_writeresponsevalid   => open,                                                                       --              (terminated)
			av_writeresponserequest  => open,                                                                       --              (terminated)
			av_writeresponsevalid    => '0'                                                                         --              (terminated)
		);

	timer_timestamp_s1_translator : component sopc_video_timer_system_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                    reset.reset
			uav_address              => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_timestamp_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_timestamp_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_timestamp_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_timestamp_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                          --              (terminated)
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_burstcount            => open,                                                                          --              (terminated)
			av_byteenable            => open,                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_debugaccess           => open,                                                                          --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	lcd_control_slave_translator : component sopc_video_lcd_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 13,
			AV_WRITE_WAIT_CYCLES           => 13,
			AV_SETUP_WAIT_CYCLES           => 13,
			AV_DATA_HOLD_CYCLES            => 13
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address              => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lcd_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lcd_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => lcd_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => lcd_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => lcd_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_beginbursttransfer    => open,                                                                         --              (terminated)
			av_burstcount            => open,                                                                         --              (terminated)
			av_byteenable            => open,                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                         --              (terminated)
			av_lock                  => open,                                                                         --              (terminated)
			av_chipselect            => open,                                                                         --              (terminated)
			av_clken                 => open,                                                                         --              (terminated)
			uav_clken                => '0',                                                                          --              (terminated)
			av_debugaccess           => open,                                                                         --              (terminated)
			av_outputenable          => open,                                                                         --              (terminated)
			uav_response             => open,                                                                         --              (terminated)
			av_response              => "00",                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                           --              (terminated)
		);

	red_leds_s1_translator : component sopc_video_red_leds_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => red_leds_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => red_leds_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => red_leds_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => red_leds_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => red_leds_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	green_leds_s1_translator : component sopc_video_red_leds_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => green_leds_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => green_leds_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => green_leds_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => green_leds_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => green_leds_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	switch_s1_translator : component sopc_video_switch_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => switch_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => switch_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => switch_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => switch_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => switch_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => switch_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                 --              (terminated)
			av_read                  => open,                                                                 --              (terminated)
			av_writedata             => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_chipselect            => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator : component sopc_video_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                                                      --                    reset.reset
			uav_address              => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                                                                --              (terminated)
			av_burstcount            => open,                                                                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                                                                --              (terminated)
			av_lock                  => open,                                                                                                                --              (terminated)
			av_clken                 => open,                                                                                                                --              (terminated)
			uav_clken                => '0',                                                                                                                 --              (terminated)
			av_debugaccess           => open,                                                                                                                --              (terminated)
			av_outputenable          => open,                                                                                                                --              (terminated)
			uav_response             => open,                                                                                                                --              (terminated)
			av_response              => "00",                                                                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                                                                  --              (terminated)
		);

	barcode_scan_0_s1_translator : component sopc_video_barcode_scan_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 8,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 1,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 1,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 1,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clock_signals_sys_clk_clk,                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address              => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => barcode_scan_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => barcode_scan_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => barcode_scan_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => barcode_scan_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => barcode_scan_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => barcode_scan_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                         --              (terminated)
			av_burstcount            => open,                                                                         --              (terminated)
			av_byteenable            => open,                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                         --              (terminated)
			av_lock                  => open,                                                                         --              (terminated)
			av_clken                 => open,                                                                         --              (terminated)
			uav_clken                => '0',                                                                          --              (terminated)
			av_debugaccess           => open,                                                                         --              (terminated)
			av_outputenable          => open,                                                                         --              (terminated)
			uav_response             => open,                                                                         --              (terminated)
			av_response              => "00",                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                           --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component sopc_video_cpu_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_BEGIN_BURST           => 87,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			PKT_BURST_TYPE_H          => 84,
			PKT_BURST_TYPE_L          => 83,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_THREAD_ID_H           => 99,
			PKT_THREAD_ID_L           => 99,
			PKT_CACHE_H               => 106,
			PKT_CACHE_L               => 103,
			PKT_DATA_SIDEBAND_H       => 86,
			PKT_DATA_SIDEBAND_L       => 86,
			PKT_QOS_H                 => 88,
			PKT_QOS_L                 => 88,
			PKT_ADDR_SIDEBAND_H       => 85,
			PKT_ADDR_SIDEBAND_L       => 85,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			ST_DATA_W                 => 109,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                          --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                             --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                              --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                           --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                             --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component sopc_video_cpu_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_BEGIN_BURST           => 87,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			PKT_BURST_TYPE_H          => 84,
			PKT_BURST_TYPE_L          => 83,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_THREAD_ID_H           => 99,
			PKT_THREAD_ID_L           => 99,
			PKT_CACHE_H               => 106,
			PKT_CACHE_L               => 103,
			PKT_DATA_SIDEBAND_H       => 86,
			PKT_DATA_SIDEBAND_L       => 86,
			PKT_QOS_H                 => 88,
			PKT_QOS_L                 => 88,
			PKT_ADDR_SIDEBAND_H       => 85,
			PKT_ADDR_SIDEBAND_L       => 85,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			ST_DATA_W                 => 109,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                   --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent : component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_BEGIN_BURST           => 60,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			PKT_BURST_TYPE_H          => 57,
			PKT_BURST_TYPE_L          => 56,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_POSTED          => 42,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			PKT_TRANS_LOCK            => 45,
			PKT_TRANS_EXCLUSIVE       => 46,
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_SRC_ID_H              => 66,
			PKT_SRC_ID_L              => 62,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 67,
			PKT_THREAD_ID_H           => 72,
			PKT_THREAD_ID_L           => 72,
			PKT_CACHE_H               => 79,
			PKT_CACHE_L               => 76,
			PKT_DATA_SIDEBAND_H       => 59,
			PKT_DATA_SIDEBAND_L       => 59,
			PKT_QOS_H                 => 61,
			PKT_QOS_L                 => 61,
			PKT_ADDR_SIDEBAND_H       => 58,
			PKT_ADDR_SIDEBAND_L       => 58,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 1,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 2,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                            --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                       -- clk_reset.reset
			av_address              => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => width_adapter_009_src_valid,                                                                          --        rp.valid
			rp_data                 => width_adapter_009_src_data,                                                                           --          .data
			rp_channel              => width_adapter_009_src_channel,                                                                        --          .channel
			rp_startofpacket        => width_adapter_009_src_startofpacket,                                                                  --          .startofpacket
			rp_endofpacket          => width_adapter_009_src_endofpacket,                                                                    --          .endofpacket
			rp_ready                => width_adapter_009_src_ready,                                                                          --          .ready
			av_response             => open,                                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                                  -- (terminated)
		);

	video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent : component sopc_video_pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_BEGIN_BURST           => 60,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			PKT_BURST_TYPE_H          => 57,
			PKT_BURST_TYPE_L          => 56,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_POSTED          => 42,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			PKT_TRANS_LOCK            => 45,
			PKT_TRANS_EXCLUSIVE       => 46,
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_SRC_ID_H              => 66,
			PKT_SRC_ID_L              => 62,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 67,
			PKT_THREAD_ID_H           => 72,
			PKT_THREAD_ID_L           => 72,
			PKT_CACHE_H               => 79,
			PKT_CACHE_L               => 76,
			PKT_DATA_SIDEBAND_H       => 59,
			PKT_DATA_SIDEBAND_L       => 59,
			PKT_QOS_H                 => 61,
			PKT_QOS_L                 => 61,
			PKT_ADDR_SIDEBAND_H       => 58,
			PKT_ADDR_SIDEBAND_L       => 58,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 17,
			AV_BURSTCOUNT_W           => 1,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 3,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                               --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			av_address              => video_dma_avalon_dma_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => video_dma_avalon_dma_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => video_dma_avalon_dma_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => width_adapter_010_src_valid,                                                             --        rp.valid
			rp_data                 => width_adapter_010_src_data,                                                              --          .data
			rp_channel              => width_adapter_010_src_channel,                                                           --          .channel
			rp_startofpacket        => width_adapter_010_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => width_adapter_010_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => width_adapter_010_src_ready,                                                             --          .ready
			av_response             => open,                                                                                    -- (terminated)
			av_writeresponserequest => '0',                                                                                     -- (terminated)
			av_writeresponsevalid   => open                                                                                     -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                          --                .channel
			rf_sink_ready           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 69,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 71,
			PKT_DEST_ID_H             => 80,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 84,
			PKT_PROTECTION_L          => 82,
			PKT_RESPONSE_STATUS_H     => 90,
			PKT_RESPONSE_STATUS_L     => 89,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 91,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                     --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                     --                .valid
			cp_data                 => burst_adapter_source0_data,                                                      --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                               --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                   --                .channel
			rf_sink_ready           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 92,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                            -- clk_reset.reset
			in_data           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                      -- (terminated)
			csr_read          => '0',                                                                       -- (terminated)
			csr_write         => '0',                                                                       -- (terminated)
			csr_readdata      => open,                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                        -- (terminated)
			almost_full_data  => open,                                                                      -- (terminated)
			almost_empty_data => open,                                                                      -- (terminated)
			in_startofpacket  => '0',                                                                       -- (terminated)
			in_endofpacket    => '0',                                                                       -- (terminated)
			out_startofpacket => open,                                                                      -- (terminated)
			out_endofpacket   => open,                                                                      -- (terminated)
			in_empty          => '0',                                                                       -- (terminated)
			out_empty         => open,                                                                      -- (terminated)
			in_error          => '0',                                                                       -- (terminated)
			out_error         => open,                                                                      -- (terminated)
			in_channel        => '0',                                                                       -- (terminated)
			out_channel       => open                                                                       -- (terminated)
		);

	pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 69,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 75,
			PKT_SRC_ID_L              => 71,
			PKT_DEST_ID_H             => 80,
			PKT_DEST_ID_L             => 76,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 84,
			PKT_PROTECTION_L          => 82,
			PKT_RESPONSE_STATUS_H     => 90,
			PKT_RESPONSE_STATUS_L     => 89,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 91,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                           --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                                     --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                                     --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                                      --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                               --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                                   --                .channel
			rf_sink_ready           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 92,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                           --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component sopc_video_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 3,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			in_data           => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                          -- (terminated)
			csr_read          => '0',                                                                                           -- (terminated)
			csr_write         => '0',                                                                                           -- (terminated)
			csr_readdata      => open,                                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                            -- (terminated)
			almost_full_data  => open,                                                                                          -- (terminated)
			almost_empty_data => open,                                                                                          -- (terminated)
			in_startofpacket  => '0',                                                                                           -- (terminated)
			in_endofpacket    => '0',                                                                                           -- (terminated)
			out_startofpacket => open,                                                                                          -- (terminated)
			out_endofpacket   => open,                                                                                          -- (terminated)
			in_empty          => '0',                                                                                           -- (terminated)
			out_empty         => open,                                                                                          -- (terminated)
			in_error          => '0',                                                                                           -- (terminated)
			out_error         => open,                                                                                          -- (terminated)
			in_channel        => '0',                                                                                           -- (terminated)
			out_channel       => open                                                                                           -- (terminated)
		);

	av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                        --       clk_reset.reset
			m0_address              => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                                         --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                                                       --                .channel
			rf_sink_ready           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                    --     (terminated)
		);

	av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                        -- clk_reset.reset
			in_data           => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                  -- (terminated)
			csr_read          => '0',                                                                                                   -- (terminated)
			csr_write         => '0',                                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                    -- (terminated)
			almost_full_data  => open,                                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                                  -- (terminated)
			in_empty          => '0',                                                                                                   -- (terminated)
			out_empty         => open,                                                                                                  -- (terminated)
			in_error          => '0',                                                                                                   -- (terminated)
			out_error         => open,                                                                                                  -- (terminated)
			in_channel        => '0',                                                                                                   -- (terminated)
			out_channel       => open                                                                                                   -- (terminated)
		);

	video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                          --       clk_reset.reset
			m0_address              => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                                           --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                                           --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                                            --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                                                     --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                                                         --                .channel
			rf_sink_ready           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                      --     (terminated)
		);

	video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                          -- clk_reset.reset
			in_data           => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                    -- (terminated)
			csr_read          => '0',                                                                                                     -- (terminated)
			csr_write         => '0',                                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                      -- (terminated)
			almost_full_data  => open,                                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                                    -- (terminated)
			in_empty          => '0',                                                                                                     -- (terminated)
			out_empty         => open,                                                                                                    -- (terminated)
			in_error          => '0',                                                                                                     -- (terminated)
			out_error         => open,                                                                                                    -- (terminated)
			in_channel        => '0',                                                                                                     -- (terminated)
			out_channel       => open                                                                                                     -- (terminated)
		);

	pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                             --       clk_reset.reset
			m0_address              => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                                            --                .channel
			rf_sink_ready           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                         --     (terminated)
		);

	pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                             -- clk_reset.reset
			in_data           => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                       -- (terminated)
			csr_read          => '0',                                                                                                        -- (terminated)
			csr_write         => '0',                                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                         -- (terminated)
			almost_full_data  => open,                                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                                       -- (terminated)
			in_empty          => '0',                                                                                                        -- (terminated)
			out_empty         => open,                                                                                                       -- (terminated)
			in_error          => '0',                                                                                                        -- (terminated)
			out_error         => open,                                                                                                       -- (terminated)
			in_channel        => '0',                                                                                                        -- (terminated)
			out_channel       => open                                                                                                        -- (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                                    --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                                 --                .channel
			rf_sink_ready           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                              --     (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                            -- (terminated)
			csr_read          => '0',                                                                                             -- (terminated)
			csr_write         => '0',                                                                                             -- (terminated)
			csr_readdata      => open,                                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                              -- (terminated)
			almost_full_data  => open,                                                                                            -- (terminated)
			almost_empty_data => open,                                                                                            -- (terminated)
			in_empty          => '0',                                                                                             -- (terminated)
			out_empty         => open,                                                                                            -- (terminated)
			in_error          => '0',                                                                                             -- (terminated)
			out_error         => open,                                                                                            -- (terminated)
			in_channel        => '0',                                                                                             -- (terminated)
			out_channel       => open                                                                                             -- (terminated)
		);

	timer_system_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                      --                .channel
			rf_sink_ready           => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                 --     (terminated)
			m0_writeresponserequest => open,                                                                                 --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                   --     (terminated)
		);

	timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                 -- (terminated)
			csr_read          => '0',                                                                                  -- (terminated)
			csr_write         => '0',                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                   -- (terminated)
			almost_full_data  => open,                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                 -- (terminated)
			in_empty          => '0',                                                                                  -- (terminated)
			out_empty         => open,                                                                                 -- (terminated)
			in_error          => '0',                                                                                  -- (terminated)
			out_error         => open,                                                                                 -- (terminated)
			in_channel        => '0',                                                                                  -- (terminated)
			out_channel       => open                                                                                  -- (terminated)
		);

	timer_timestamp_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src10_ready,                                                          --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src10_valid,                                                          --                .valid
			cp_data                 => cmd_xbar_demux_001_src10_data,                                                           --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src10_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src10_endofpacket,                                                    --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src10_channel,                                                        --                .channel
			rf_sink_ready           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                      --     (terminated)
		);

	timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                    -- (terminated)
			csr_read          => '0',                                                                                     -- (terminated)
			csr_write         => '0',                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                      -- (terminated)
			almost_full_data  => open,                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                    -- (terminated)
			in_empty          => '0',                                                                                     -- (terminated)
			out_empty         => open,                                                                                    -- (terminated)
			in_error          => '0',                                                                                     -- (terminated)
			out_error         => open,                                                                                    -- (terminated)
			in_channel        => '0',                                                                                     -- (terminated)
			out_channel       => open                                                                                     -- (terminated)
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src11_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src11_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_demux_001_src11_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src11_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src11_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src11_channel,                                                       --                .channel
			rf_sink_ready           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                     --     (terminated)
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                   -- (terminated)
			csr_read          => '0',                                                                                    -- (terminated)
			csr_write         => '0',                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                     -- (terminated)
			almost_full_data  => open,                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                   -- (terminated)
			in_empty          => '0',                                                                                    -- (terminated)
			out_empty         => open,                                                                                   -- (terminated)
			in_error          => '0',                                                                                    -- (terminated)
			out_error         => open,                                                                                   -- (terminated)
			in_channel        => '0',                                                                                    -- (terminated)
			out_channel       => open                                                                                    -- (terminated)
		);

	red_leds_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => red_leds_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src12_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src12_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src12_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src12_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src12_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src12_channel,                                                 --                .channel
			rf_sink_ready           => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => red_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => red_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => red_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	green_leds_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src13_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src13_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src13_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src13_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src13_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src13_channel,                                                   --                .channel
			rf_sink_ready           => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	switch_s1_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => switch_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => switch_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => switch_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => switch_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => switch_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => switch_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => switch_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src14_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src14_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src14_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src14_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src14_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src14_channel,                                               --                .channel
			rf_sink_ready           => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 87,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 93,
			PKT_SRC_ID_L              => 89,
			PKT_DEST_ID_H             => 98,
			PKT_DEST_ID_L             => 94,
			PKT_BURSTWRAP_H           => 79,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 102,
			PKT_PROTECTION_L          => 100,
			PKT_RESPONSE_STATUS_H     => 108,
			PKT_RESPONSE_STATUS_L     => 107,
			PKT_BURST_SIZE_H          => 82,
			PKT_BURST_SIZE_L          => 80,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 109,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                                                --       clk_reset.reset
			m0_address              => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src15_ready,                                                                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src15_valid,                                                                                                --                .valid
			cp_data                 => cmd_xbar_demux_001_src15_data,                                                                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src15_startofpacket,                                                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src15_endofpacket,                                                                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src15_channel,                                                                                              --                .channel
			rf_sink_ready           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                                            --     (terminated)
		);

	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 110,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                                                -- clk_reset.reset
			in_data           => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                                          -- (terminated)
			csr_read          => '0',                                                                                                                           -- (terminated)
			csr_write         => '0',                                                                                                                           -- (terminated)
			csr_readdata      => open,                                                                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                                            -- (terminated)
			almost_full_data  => open,                                                                                                                          -- (terminated)
			almost_empty_data => open,                                                                                                                          -- (terminated)
			in_empty          => '0',                                                                                                                           -- (terminated)
			out_empty         => open,                                                                                                                          -- (terminated)
			in_error          => '0',                                                                                                                           -- (terminated)
			out_error         => open,                                                                                                                          -- (terminated)
			in_channel        => '0',                                                                                                                           -- (terminated)
			out_channel       => open                                                                                                                           -- (terminated)
		);

	barcode_scan_0_s1_translator_avalon_universal_slave_0_agent : component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 60,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_POSTED          => 42,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			PKT_TRANS_LOCK            => 45,
			PKT_SRC_ID_H              => 66,
			PKT_SRC_ID_L              => 62,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 67,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			ST_CHANNEL_W              => 17,
			ST_DATA_W                 => 82,
			AVS_BURSTCOUNT_W          => 1,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clock_signals_sys_clk_clk,                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_002_source0_ready,                                                        --              cp.ready
			cp_valid                => burst_adapter_002_source0_valid,                                                        --                .valid
			cp_data                 => burst_adapter_002_source0_data,                                                         --                .data
			cp_startofpacket        => burst_adapter_002_source0_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => burst_adapter_002_source0_endofpacket,                                                  --                .endofpacket
			cp_channel              => burst_adapter_002_source0_channel,                                                      --                .channel
			rf_sink_ready           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                     --     (terminated)
		);

	barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_video_barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 83,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clock_signals_sys_clk_clk,                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                   -- (terminated)
			csr_read          => '0',                                                                                    -- (terminated)
			csr_write         => '0',                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                     -- (terminated)
			almost_full_data  => open,                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                   -- (terminated)
			in_empty          => '0',                                                                                    -- (terminated)
			out_empty         => open,                                                                                   -- (terminated)
			in_error          => '0',                                                                                    -- (terminated)
			out_error         => open,                                                                                   -- (terminated)
			in_channel        => '0',                                                                                    -- (terminated)
			out_channel       => open                                                                                    -- (terminated)
		);

	addr_router : component SOPC_Video_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component SOPC_Video_addr_router_001
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                   --       src.ready
			src_valid          => addr_router_001_src_valid,                                                   --          .valid
			src_data           => addr_router_001_src_data,                                                    --          .data
			src_channel        => addr_router_001_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                              --          .endofpacket
		);

	addr_router_002 : component SOPC_Video_addr_router_002
		port map (
			sink_ready         => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                       -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                                                            --       src.ready
			src_valid          => addr_router_002_src_valid,                                                                            --          .valid
			src_data           => addr_router_002_src_data,                                                                             --          .data
			src_channel        => addr_router_002_src_channel,                                                                          --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                                                    --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                                                       --          .endofpacket
		);

	addr_router_003 : component SOPC_Video_addr_router_002
		port map (
			sink_ready         => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => addr_router_003_src_ready,                                                               --       src.ready
			src_valid          => addr_router_003_src_valid,                                                               --          .valid
			src_data           => addr_router_003_src_data,                                                                --          .data
			src_channel        => addr_router_003_src_channel,                                                             --          .channel
			src_startofpacket  => addr_router_003_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => addr_router_003_src_endofpacket                                                          --          .endofpacket
		);

	id_router : component SOPC_Video_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component SOPC_Video_id_router
		port map (
			sink_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                     --       src.ready
			src_valid          => id_router_001_src_valid,                                                     --          .valid
			src_data           => id_router_001_src_data,                                                      --          .data
			src_channel        => id_router_001_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                --          .endofpacket
		);

	id_router_002 : component SOPC_Video_id_router_002
		port map (
			sink_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                               --       src.ready
			src_valid          => id_router_002_src_valid,                                               --          .valid
			src_data           => id_router_002_src_data,                                                --          .data
			src_channel        => id_router_002_src_channel,                                             --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                          --          .endofpacket
		);

	id_router_003 : component SOPC_Video_id_router_003
		port map (
			sink_ready         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                                   --       src.ready
			src_valid          => id_router_003_src_valid,                                                                   --          .valid
			src_data           => id_router_003_src_data,                                                                    --          .data
			src_channel        => id_router_003_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                              --          .endofpacket
		);

	id_router_004 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                     --       src.ready
			src_valid          => id_router_004_src_valid,                                                                     --          .valid
			src_data           => id_router_004_src_data,                                                                      --          .data
			src_channel        => id_router_004_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                                --          .endofpacket
		);

	id_router_005 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                                       --       src.ready
			src_valid          => id_router_005_src_valid,                                                                       --          .valid
			src_data           => id_router_005_src_data,                                                                        --          .data
			src_channel        => id_router_005_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                                  --          .endofpacket
		);

	id_router_006 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                          --       src.ready
			src_valid          => id_router_006_src_valid,                                                                          --          .valid
			src_data           => id_router_006_src_data,                                                                           --          .data
			src_channel        => id_router_006_src_channel,                                                                        --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                                  --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                                     --          .endofpacket
		);

	id_router_007 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                                  --       src.ready
			src_valid          => id_router_007_src_valid,                                                                  --          .valid
			src_data           => id_router_007_src_data,                                                                   --          .data
			src_channel        => id_router_007_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                             --          .endofpacket
		);

	id_router_008 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                               --       src.ready
			src_valid          => id_router_008_src_valid,                                                               --          .valid
			src_data           => id_router_008_src_data,                                                                --          .data
			src_channel        => id_router_008_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                          --          .endofpacket
		);

	id_router_009 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                    --       src.ready
			src_valid          => id_router_009_src_valid,                                                    --          .valid
			src_data           => id_router_009_src_data,                                                     --          .data
			src_channel        => id_router_009_src_channel,                                                  --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                            --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                               --          .endofpacket
		);

	id_router_010 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                       --       src.ready
			src_valid          => id_router_010_src_valid,                                                       --          .valid
			src_data           => id_router_010_src_data,                                                        --          .data
			src_channel        => id_router_010_src_channel,                                                     --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                                  --          .endofpacket
		);

	id_router_011 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                      --       src.ready
			src_valid          => id_router_011_src_valid,                                                      --          .valid
			src_data           => id_router_011_src_data,                                                       --          .data
			src_channel        => id_router_011_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                                 --          .endofpacket
		);

	id_router_012 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => red_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                --       src.ready
			src_valid          => id_router_012_src_valid,                                                --          .valid
			src_data           => id_router_012_src_data,                                                 --          .data
			src_channel        => id_router_012_src_channel,                                              --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                           --          .endofpacket
		);

	id_router_013 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                  --       src.ready
			src_valid          => id_router_013_src_valid,                                                  --          .valid
			src_data           => id_router_013_src_data,                                                   --          .data
			src_channel        => id_router_013_src_channel,                                                --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                             --          .endofpacket
		);

	id_router_014 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => switch_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => switch_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => switch_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                              --       src.ready
			src_valid          => id_router_014_src_valid,                                              --          .valid
			src_data           => id_router_014_src_data,                                               --          .data
			src_channel        => id_router_014_src_channel,                                            --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                         --          .endofpacket
		);

	id_router_015 : component SOPC_Video_id_router_004
		port map (
			sink_ready         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                                      -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                                                                             --       src.ready
			src_valid          => id_router_015_src_valid,                                                                                             --          .valid
			src_data           => id_router_015_src_data,                                                                                              --          .data
			src_channel        => id_router_015_src_channel,                                                                                           --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                                                                     --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                                                                        --          .endofpacket
		);

	id_router_016 : component SOPC_Video_id_router_016
		port map (
			sink_ready         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => barcode_scan_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clock_signals_sys_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                                      --       src.ready
			src_valid          => id_router_016_src_valid,                                                      --          .valid
			src_data           => id_router_016_src_data,                                                       --          .data
			src_channel        => id_router_016_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                                 --          .endofpacket
		);

	burst_adapter : component sopc_video_burst_adapter
		generic map (
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 69,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			PKT_BURST_TYPE_H          => 66,
			PKT_BURST_TYPE_L          => 65,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 91,
			ST_CHANNEL_W              => 17,
			OUT_BYTE_CNT_H            => 57,
			OUT_BURSTWRAP_H           => 61,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clock_signals_sys_clk_clk,           --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_002_src_valid,          --     sink0.valid
			sink0_data            => cmd_xbar_mux_002_src_data,           --          .data
			sink0_channel         => cmd_xbar_mux_002_src_channel,        --          .channel
			sink0_startofpacket   => cmd_xbar_mux_002_src_startofpacket,  --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_002_src_endofpacket,    --          .endofpacket
			sink0_ready           => cmd_xbar_mux_002_src_ready,          --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component sopc_video_burst_adapter
		generic map (
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 69,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 64,
			PKT_BURST_SIZE_L          => 62,
			PKT_BURST_TYPE_H          => 66,
			PKT_BURST_TYPE_L          => 65,
			PKT_BURSTWRAP_H           => 61,
			PKT_BURSTWRAP_L           => 59,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 91,
			ST_CHANNEL_W              => 17,
			OUT_BYTE_CNT_H            => 57,
			OUT_BURSTWRAP_H           => 61,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 7,
			BURSTWRAP_CONST_VALUE     => 7
		)
		port map (
			clk                   => clock_signals_sys_clk_clk,               --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_003_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_003_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_003_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_003_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_003_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_003_src_ready,              --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	burst_adapter_002 : component sopc_video_burst_adapter_002
		generic map (
			PKT_ADDR_H                => 40,
			PKT_ADDR_L                => 9,
			PKT_BEGIN_BURST           => 60,
			PKT_BYTE_CNT_H            => 49,
			PKT_BYTE_CNT_L            => 47,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_BURST_SIZE_H          => 55,
			PKT_BURST_SIZE_L          => 53,
			PKT_BURST_TYPE_H          => 57,
			PKT_BURST_TYPE_L          => 56,
			PKT_BURSTWRAP_H           => 52,
			PKT_BURSTWRAP_L           => 50,
			PKT_TRANS_COMPRESSED_READ => 41,
			PKT_TRANS_WRITE           => 43,
			PKT_TRANS_READ            => 44,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 17,
			OUT_BYTE_CNT_H            => 47,
			OUT_BURSTWRAP_H           => 52,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 7,
			BURSTWRAP_CONST_VALUE     => 7
		)
		port map (
			clk                   => clock_signals_sys_clk_clk,               --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => width_adapter_003_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_003_src_data,              --          .data
			sink0_channel         => width_adapter_003_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_003_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_003_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_003_src_ready,             --          .ready
			source0_valid         => burst_adapter_002_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_002_source0_data,          --          .data
			source0_channel       => burst_adapter_002_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_002_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_002_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_002_source0_ready          --          .ready
		);

	rst_controller : component sopc_video_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 4,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => reset_n_ports_inv,                           -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,           -- reset_in1.reset
			reset_in2  => clock_signals_sys_clk_reset_reset_ports_inv, -- reset_in2.reset
			reset_in3  => rst_controller_003_reset_out_reset,          -- reset_in3.reset
			clk        => clock_signals_sys_clk_clk,                   --       clk.clk
			reset_out  => rst_controller_reset_out_reset,              -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req,          --          .reset_req
			reset_in4  => '0',                                         -- (terminated)
			reset_in5  => '0',                                         -- (terminated)
			reset_in6  => '0',                                         -- (terminated)
			reset_in7  => '0',                                         -- (terminated)
			reset_in8  => '0',                                         -- (terminated)
			reset_in9  => '0',                                         -- (terminated)
			reset_in10 => '0',                                         -- (terminated)
			reset_in11 => '0',                                         -- (terminated)
			reset_in12 => '0',                                         -- (terminated)
			reset_in13 => '0',                                         -- (terminated)
			reset_in14 => '0',                                         -- (terminated)
			reset_in15 => '0'                                          -- (terminated)
		);

	rst_controller_001 : component sopc_video_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 4,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                           -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,           -- reset_in1.reset
			reset_in2  => clock_signals_sys_clk_reset_reset_ports_inv, -- reset_in2.reset
			reset_in3  => rst_controller_003_reset_out_reset,          -- reset_in3.reset
			clk        => clock_signals_vga_clk_clk,                   --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,          -- reset_out.reset
			reset_req  => open,                                        -- (terminated)
			reset_in4  => '0',                                         -- (terminated)
			reset_in5  => '0',                                         -- (terminated)
			reset_in6  => '0',                                         -- (terminated)
			reset_in7  => '0',                                         -- (terminated)
			reset_in8  => '0',                                         -- (terminated)
			reset_in9  => '0',                                         -- (terminated)
			reset_in10 => '0',                                         -- (terminated)
			reset_in11 => '0',                                         -- (terminated)
			reset_in12 => '0',                                         -- (terminated)
			reset_in13 => '0',                                         -- (terminated)
			reset_in14 => '0',                                         -- (terminated)
			reset_in15 => '0'                                          -- (terminated)
		);

	rst_controller_002 : component sopc_video_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 4,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                           -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,           -- reset_in1.reset
			reset_in2  => clock_signals_sys_clk_reset_reset_ports_inv, -- reset_in2.reset
			reset_in3  => rst_controller_003_reset_out_reset,          -- reset_in3.reset
			clk        => clk_0,                                       --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset,          -- reset_out.reset
			reset_req  => open,                                        -- (terminated)
			reset_in4  => '0',                                         -- (terminated)
			reset_in5  => '0',                                         -- (terminated)
			reset_in6  => '0',                                         -- (terminated)
			reset_in7  => '0',                                         -- (terminated)
			reset_in8  => '0',                                         -- (terminated)
			reset_in9  => '0',                                         -- (terminated)
			reset_in10 => '0',                                         -- (terminated)
			reset_in11 => '0',                                         -- (terminated)
			reset_in12 => '0',                                         -- (terminated)
			reset_in13 => '0',                                         -- (terminated)
			reset_in14 => '0',                                         -- (terminated)
			reset_in15 => '0'                                          -- (terminated)
		);

	rst_controller_003 : component sopc_video_rst_controller_003
		generic map (
			NUM_RESET_INPUTS        => 3,
			OUTPUT_RESET_SYNC_EDGES => "none",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                           -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset,           -- reset_in1.reset
			reset_in2  => clock_signals_sys_clk_reset_reset_ports_inv, -- reset_in2.reset
			clk        => open,                                        --       clk.clk
			reset_out  => rst_controller_003_reset_out_reset,          -- reset_out.reset
			reset_req  => open,                                        -- (terminated)
			reset_in3  => '0',                                         -- (terminated)
			reset_in4  => '0',                                         -- (terminated)
			reset_in5  => '0',                                         -- (terminated)
			reset_in6  => '0',                                         -- (terminated)
			reset_in7  => '0',                                         -- (terminated)
			reset_in8  => '0',                                         -- (terminated)
			reset_in9  => '0',                                         -- (terminated)
			reset_in10 => '0',                                         -- (terminated)
			reset_in11 => '0',                                         -- (terminated)
			reset_in12 => '0',                                         -- (terminated)
			reset_in13 => '0',                                         -- (terminated)
			reset_in14 => '0',                                         -- (terminated)
			reset_in15 => '0'                                          -- (terminated)
		);

	cmd_xbar_demux : component SOPC_Video_cmd_xbar_demux
		port map (
			clk                => clock_signals_sys_clk_clk,         --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component SOPC_Video_cmd_xbar_demux_001
		port map (
			clk                 => clock_signals_sys_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			sink_ready          => addr_router_001_src_ready,              --      sink.ready
			sink_channel        => addr_router_001_src_channel,            --          .channel
			sink_data           => addr_router_001_src_data,               --          .data
			sink_startofpacket  => addr_router_001_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_001_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_001_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket,   --          .endofpacket
			src14_ready         => cmd_xbar_demux_001_src14_ready,         --     src14.ready
			src14_valid         => cmd_xbar_demux_001_src14_valid,         --          .valid
			src14_data          => cmd_xbar_demux_001_src14_data,          --          .data
			src14_channel       => cmd_xbar_demux_001_src14_channel,       --          .channel
			src14_startofpacket => cmd_xbar_demux_001_src14_startofpacket, --          .startofpacket
			src14_endofpacket   => cmd_xbar_demux_001_src14_endofpacket,   --          .endofpacket
			src15_ready         => cmd_xbar_demux_001_src15_ready,         --     src15.ready
			src15_valid         => cmd_xbar_demux_001_src15_valid,         --          .valid
			src15_data          => cmd_xbar_demux_001_src15_data,          --          .data
			src15_channel       => cmd_xbar_demux_001_src15_channel,       --          .channel
			src15_startofpacket => cmd_xbar_demux_001_src15_startofpacket, --          .startofpacket
			src15_endofpacket   => cmd_xbar_demux_001_src15_endofpacket,   --          .endofpacket
			src16_ready         => cmd_xbar_demux_001_src16_ready,         --     src16.ready
			src16_valid         => cmd_xbar_demux_001_src16_valid,         --          .valid
			src16_data          => cmd_xbar_demux_001_src16_data,          --          .data
			src16_channel       => cmd_xbar_demux_001_src16_channel,       --          .channel
			src16_startofpacket => cmd_xbar_demux_001_src16_startofpacket, --          .startofpacket
			src16_endofpacket   => cmd_xbar_demux_001_src16_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_002 : component SOPC_Video_cmd_xbar_demux_002
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_002_src_ready,             --      sink.ready
			sink_channel       => addr_router_002_src_channel,           --          .channel
			sink_data          => addr_router_002_src_data,              --          .data
			sink_startofpacket => addr_router_002_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_002_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_002_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_002_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_003 : component SOPC_Video_cmd_xbar_demux_002
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_003_src_ready,             --      sink.ready
			sink_channel       => addr_router_003_src_channel,           --          .channel
			sink_data          => addr_router_003_src_data,              --          .data
			sink_startofpacket => addr_router_003_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_003_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_003_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_003_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component SOPC_Video_cmd_xbar_mux
		port map (
			clk                 => clock_signals_sys_clk_clk,             --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component SOPC_Video_cmd_xbar_mux
		port map (
			clk                 => clock_signals_sys_clk_clk,             --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component SOPC_Video_cmd_xbar_mux_002
		port map (
			clk                 => clock_signals_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,      -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,          --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,          --          .valid
			src_data            => cmd_xbar_mux_002_src_data,           --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,        --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,  --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,    --          .endofpacket
			sink0_ready         => width_adapter_src_ready,             --     sink0.ready
			sink0_valid         => width_adapter_src_valid,             --          .valid
			sink0_channel       => width_adapter_src_channel,           --          .channel
			sink0_data          => width_adapter_src_data,              --          .data
			sink0_startofpacket => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket   => width_adapter_src_endofpacket,       --          .endofpacket
			sink1_ready         => width_adapter_001_src_ready,         --     sink1.ready
			sink1_valid         => width_adapter_001_src_valid,         --          .valid
			sink1_channel       => width_adapter_001_src_channel,       --          .channel
			sink1_data          => width_adapter_001_src_data,          --          .data
			sink1_startofpacket => width_adapter_001_src_startofpacket, --          .startofpacket
			sink1_endofpacket   => width_adapter_001_src_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component SOPC_Video_cmd_xbar_mux_003
		port map (
			clk                 => clock_signals_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,      -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,          --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,          --          .valid
			src_data            => cmd_xbar_mux_003_src_data,           --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,        --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,  --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,    --          .endofpacket
			sink0_ready         => width_adapter_002_src_ready,         --     sink0.ready
			sink0_valid         => width_adapter_002_src_valid,         --          .valid
			sink0_channel       => width_adapter_002_src_channel,       --          .channel
			sink0_data          => width_adapter_002_src_data,          --          .data
			sink0_startofpacket => width_adapter_002_src_startofpacket, --          .startofpacket
			sink0_endofpacket   => width_adapter_002_src_endofpacket,   --          .endofpacket
			sink1_ready         => width_adapter_004_src_ready,         --     sink1.ready
			sink1_valid         => width_adapter_004_src_valid,         --          .valid
			sink1_channel       => width_adapter_004_src_channel,       --          .channel
			sink1_data          => width_adapter_004_src_data,          --          .data
			sink1_startofpacket => width_adapter_004_src_startofpacket, --          .startofpacket
			sink1_endofpacket   => width_adapter_004_src_endofpacket,   --          .endofpacket
			sink2_ready         => width_adapter_005_src_ready,         --     sink2.ready
			sink2_valid         => width_adapter_005_src_valid,         --          .valid
			sink2_channel       => width_adapter_005_src_channel,       --          .channel
			sink2_data          => width_adapter_005_src_data,          --          .data
			sink2_startofpacket => width_adapter_005_src_startofpacket, --          .startofpacket
			sink2_endofpacket   => width_adapter_005_src_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component SOPC_Video_rsp_xbar_demux
		port map (
			clk                => clock_signals_sys_clk_clk,         --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component SOPC_Video_rsp_xbar_demux
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component SOPC_Video_rsp_xbar_demux_002
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component SOPC_Video_rsp_xbar_demux_003
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_003_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_003_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_003_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_003_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_003_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_003_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component SOPC_Video_rsp_xbar_demux_004
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component SOPC_Video_cmd_xbar_demux_002
		port map (
			clk                => clock_signals_sys_clk_clk,             --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component SOPC_Video_rsp_xbar_mux
		port map (
			clk                 => clock_signals_sys_clk_clk,             --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => width_adapter_006_src_ready,           --     sink2.ready
			sink2_valid         => width_adapter_006_src_valid,           --          .valid
			sink2_channel       => width_adapter_006_src_channel,         --          .channel
			sink2_data          => width_adapter_006_src_data,            --          .data
			sink2_startofpacket => width_adapter_006_src_startofpacket,   --          .startofpacket
			sink2_endofpacket   => width_adapter_006_src_endofpacket      --          .endofpacket
		);

	rsp_xbar_mux_001 : component SOPC_Video_rsp_xbar_mux_001
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => width_adapter_007_src_ready,           --     sink2.ready
			sink2_valid          => width_adapter_007_src_valid,           --          .valid
			sink2_channel        => width_adapter_007_src_channel,         --          .channel
			sink2_data           => width_adapter_007_src_data,            --          .data
			sink2_startofpacket  => width_adapter_007_src_startofpacket,   --          .startofpacket
			sink2_endofpacket    => width_adapter_007_src_endofpacket,     --          .endofpacket
			sink3_ready          => width_adapter_008_src_ready,           --     sink3.ready
			sink3_valid          => width_adapter_008_src_valid,           --          .valid
			sink3_channel        => width_adapter_008_src_channel,         --          .channel
			sink3_data           => width_adapter_008_src_data,            --          .data
			sink3_startofpacket  => width_adapter_008_src_startofpacket,   --          .startofpacket
			sink3_endofpacket    => width_adapter_008_src_endofpacket,     --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src0_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink16_ready         => width_adapter_011_src_ready,           --    sink16.ready
			sink16_valid         => width_adapter_011_src_valid,           --          .valid
			sink16_channel       => width_adapter_011_src_channel,         --          .channel
			sink16_data          => width_adapter_011_src_data,            --          .data
			sink16_startofpacket => width_adapter_011_src_startofpacket,   --          .startofpacket
			sink16_endofpacket   => width_adapter_011_src_endofpacket      --          .endofpacket
		);

	width_adapter : component sopc_video_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,         --       clk.clk
			reset                => rst_controller_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src2_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_src2_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_src2_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src2_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_src2_ready,         --          .ready
			in_data              => cmd_xbar_demux_src2_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_src_data,            --          .data
			out_channel          => width_adapter_src_channel,         --          .channel
			out_valid            => width_adapter_src_valid,           --          .valid
			out_ready            => width_adapter_src_ready,           --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                              -- (terminated)
		);

	width_adapter_001 : component sopc_video_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src2_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src2_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src2_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src2_data,          --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_001_src_data,            --          .data
			out_channel          => width_adapter_001_src_channel,         --          .channel
			out_valid            => width_adapter_001_src_valid,           --          .valid
			out_ready            => width_adapter_001_src_ready,           --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_002 : component sopc_video_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src3_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src3_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src3_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src3_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src3_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_002_src_data,            --          .data
			out_channel          => width_adapter_002_src_channel,         --          .channel
			out_valid            => width_adapter_002_src_valid,           --          .valid
			out_ready            => width_adapter_002_src_ready,           --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_003 : component sopc_video_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 76,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 79,
			IN_PKT_BURSTWRAP_L            => 77,
			IN_PKT_BURST_SIZE_H           => 82,
			IN_PKT_BURST_SIZE_L           => 80,
			IN_PKT_RESPONSE_STATUS_H      => 108,
			IN_PKT_RESPONSE_STATUS_L      => 107,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 84,
			IN_PKT_BURST_TYPE_L           => 83,
			IN_ST_DATA_W                  => 109,
			OUT_PKT_ADDR_H                => 40,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 49,
			OUT_PKT_BYTE_CNT_L            => 47,
			OUT_PKT_TRANS_COMPRESSED_READ => 41,
			OUT_PKT_BURST_SIZE_H          => 55,
			OUT_PKT_BURST_SIZE_L          => 53,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 46,
			OUT_PKT_BURST_TYPE_H          => 57,
			OUT_PKT_BURST_TYPE_L          => 56,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,              --       clk.clk
			reset                => rst_controller_reset_out_reset,         -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src16_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src16_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src16_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src16_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src16_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src16_data,          --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_003_src_data,             --          .data
			out_channel          => width_adapter_003_src_channel,          --          .channel
			out_valid            => width_adapter_003_src_valid,            --          .valid
			out_ready            => width_adapter_003_src_ready,            --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                                   -- (terminated)
		);

	width_adapter_004 : component sopc_video_width_adapter_004
		generic map (
			IN_PKT_ADDR_H                 => 40,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 49,
			IN_PKT_BYTE_CNT_L             => 47,
			IN_PKT_TRANS_COMPRESSED_READ  => 41,
			IN_PKT_BURSTWRAP_H            => 52,
			IN_PKT_BURSTWRAP_L            => 50,
			IN_PKT_BURST_SIZE_H           => 55,
			IN_PKT_BURST_SIZE_L           => 53,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 46,
			IN_PKT_BURST_TYPE_H           => 57,
			IN_PKT_BURST_TYPE_L           => 56,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_002_src0_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_002_src0_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_002_src0_ready,         --          .ready
			in_data              => cmd_xbar_demux_002_src0_data,          --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_004_src_data,            --          .data
			out_channel          => width_adapter_004_src_channel,         --          .channel
			out_valid            => width_adapter_004_src_valid,           --          .valid
			out_ready            => width_adapter_004_src_ready,           --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_005 : component sopc_video_width_adapter_004
		generic map (
			IN_PKT_ADDR_H                 => 40,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 49,
			IN_PKT_BYTE_CNT_L             => 47,
			IN_PKT_TRANS_COMPRESSED_READ  => 41,
			IN_PKT_BURSTWRAP_H            => 52,
			IN_PKT_BURSTWRAP_L            => 50,
			IN_PKT_BURST_SIZE_H           => 55,
			IN_PKT_BURST_SIZE_L           => 53,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 46,
			IN_PKT_BURST_TYPE_H           => 57,
			IN_PKT_BURST_TYPE_L           => 56,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 58,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 64,
			OUT_PKT_BURST_SIZE_L          => 62,
			OUT_PKT_RESPONSE_STATUS_H     => 90,
			OUT_PKT_RESPONSE_STATUS_L     => 89,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 66,
			OUT_PKT_BURST_TYPE_L          => 65,
			OUT_ST_DATA_W                 => 91,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_003_src0_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_003_src0_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_003_src0_ready,         --          .ready
			in_data              => cmd_xbar_demux_003_src0_data,          --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_005_src_data,            --          .data
			out_channel          => width_adapter_005_src_channel,         --          .channel
			out_valid            => width_adapter_005_src_valid,           --          .valid
			out_ready            => width_adapter_005_src_ready,           --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_006 : component sopc_video_width_adapter_006
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_002_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_002_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_002_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_002_src0_data,          --          .data
			out_endofpacket      => width_adapter_006_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_006_src_data,            --          .data
			out_channel          => width_adapter_006_src_channel,         --          .channel
			out_valid            => width_adapter_006_src_valid,           --          .valid
			out_ready            => width_adapter_006_src_ready,           --          .ready
			out_startofpacket    => width_adapter_006_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_007 : component sopc_video_width_adapter_006
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_002_src1_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_002_src1_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_002_src1_ready,         --          .ready
			in_data              => rsp_xbar_demux_002_src1_data,          --          .data
			out_endofpacket      => width_adapter_007_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_007_src_data,            --          .data
			out_channel          => width_adapter_007_src_channel,         --          .channel
			out_valid            => width_adapter_007_src_valid,           --          .valid
			out_ready            => width_adapter_007_src_ready,           --          .ready
			out_startofpacket    => width_adapter_007_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_008 : component sopc_video_width_adapter_006
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_003_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_003_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_003_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_003_src0_data,          --          .data
			out_endofpacket      => width_adapter_008_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_008_src_data,            --          .data
			out_channel          => width_adapter_008_src_channel,         --          .channel
			out_valid            => width_adapter_008_src_valid,           --          .valid
			out_ready            => width_adapter_008_src_ready,           --          .ready
			out_startofpacket    => width_adapter_008_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_009 : component sopc_video_width_adapter_009
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 40,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 49,
			OUT_PKT_BYTE_CNT_L            => 47,
			OUT_PKT_TRANS_COMPRESSED_READ => 41,
			OUT_PKT_BURST_SIZE_H          => 55,
			OUT_PKT_BURST_SIZE_L          => 53,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 46,
			OUT_PKT_BURST_TYPE_H          => 57,
			OUT_PKT_BURST_TYPE_L          => 56,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_003_src1_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_003_src1_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_003_src1_ready,         --          .ready
			in_data              => rsp_xbar_demux_003_src1_data,          --          .data
			out_endofpacket      => width_adapter_009_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_009_src_data,            --          .data
			out_channel          => width_adapter_009_src_channel,         --          .channel
			out_valid            => width_adapter_009_src_valid,           --          .valid
			out_ready            => width_adapter_009_src_ready,           --          .ready
			out_startofpacket    => width_adapter_009_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_010 : component sopc_video_width_adapter_009
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 58,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 61,
			IN_PKT_BURSTWRAP_L            => 59,
			IN_PKT_BURST_SIZE_H           => 64,
			IN_PKT_BURST_SIZE_L           => 62,
			IN_PKT_RESPONSE_STATUS_H      => 90,
			IN_PKT_RESPONSE_STATUS_L      => 89,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 66,
			IN_PKT_BURST_TYPE_L           => 65,
			IN_ST_DATA_W                  => 91,
			OUT_PKT_ADDR_H                => 40,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 49,
			OUT_PKT_BYTE_CNT_L            => 47,
			OUT_PKT_TRANS_COMPRESSED_READ => 41,
			OUT_PKT_BURST_SIZE_H          => 55,
			OUT_PKT_BURST_SIZE_L          => 53,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 46,
			OUT_PKT_BURST_TYPE_H          => 57,
			OUT_PKT_BURST_TYPE_L          => 56,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_003_src2_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_003_src2_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_003_src2_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_003_src2_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_003_src2_ready,         --          .ready
			in_data              => rsp_xbar_demux_003_src2_data,          --          .data
			out_endofpacket      => width_adapter_010_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_010_src_data,            --          .data
			out_channel          => width_adapter_010_src_channel,         --          .channel
			out_valid            => width_adapter_010_src_valid,           --          .valid
			out_ready            => width_adapter_010_src_ready,           --          .ready
			out_startofpacket    => width_adapter_010_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_011 : component sopc_video_width_adapter_011
		generic map (
			IN_PKT_ADDR_H                 => 40,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 49,
			IN_PKT_BYTE_CNT_L             => 47,
			IN_PKT_TRANS_COMPRESSED_READ  => 41,
			IN_PKT_BURSTWRAP_H            => 52,
			IN_PKT_BURSTWRAP_L            => 50,
			IN_PKT_BURST_SIZE_H           => 55,
			IN_PKT_BURST_SIZE_L           => 53,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 46,
			IN_PKT_BURST_TYPE_H           => 57,
			IN_PKT_BURST_TYPE_L           => 56,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 76,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 82,
			OUT_PKT_BURST_SIZE_L          => 80,
			OUT_PKT_RESPONSE_STATUS_H     => 108,
			OUT_PKT_RESPONSE_STATUS_L     => 107,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 84,
			OUT_PKT_BURST_TYPE_L          => 83,
			OUT_ST_DATA_W                 => 109,
			ST_CHANNEL_W                  => 17,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clock_signals_sys_clk_clk,             --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_016_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_016_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_016_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_016_src0_data,          --          .data
			out_endofpacket      => width_adapter_011_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_011_src_data,            --          .data
			out_channel          => width_adapter_011_src_channel,         --          .channel
			out_valid            => width_adapter_011_src_valid,           --          .valid
			out_ready            => width_adapter_011_src_ready,           --          .ready
			out_startofpacket    => width_adapter_011_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	irq_mapper : component SOPC_Video_irq_mapper
		port map (
			clk           => clock_signals_sys_clk_clk,      --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	reset_n_ports_inv <= not reset_n;

	sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_write;

	sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_read;

	sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_byteenable;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	timer_system_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_system_s1_translator_avalon_anti_slave_0_write;

	timer_timestamp_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_timestamp_s1_translator_avalon_anti_slave_0_write;

	red_leds_s1_translator_avalon_anti_slave_0_write_ports_inv <= not red_leds_s1_translator_avalon_anti_slave_0_write;

	green_leds_s1_translator_avalon_anti_slave_0_write_ports_inv <= not green_leds_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	clock_signals_sys_clk_reset_reset_ports_inv <= not clock_signals_sys_clk_reset_reset;

	vga_clk <= clock_signals_vga_clk_clk;

end architecture rtl; -- of SOPC_Video
